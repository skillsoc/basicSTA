module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire net15;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire net16;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire net364;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire net2;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire net348;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire net321;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire net299;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire net14;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10493_;
 wire net17;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire net358;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire net278;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire net359;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire net292;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire net18;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire net313;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire clk_i_regs;
 wire \alu_adder_result_ex[0] ;
 wire \alu_adder_result_ex[10] ;
 wire \alu_adder_result_ex[11] ;
 wire \alu_adder_result_ex[12] ;
 wire \alu_adder_result_ex[13] ;
 wire \alu_adder_result_ex[14] ;
 wire \alu_adder_result_ex[15] ;
 wire \alu_adder_result_ex[16] ;
 wire \alu_adder_result_ex[17] ;
 wire \alu_adder_result_ex[18] ;
 wire \alu_adder_result_ex[19] ;
 wire \alu_adder_result_ex[1] ;
 wire \alu_adder_result_ex[20] ;
 wire \alu_adder_result_ex[21] ;
 wire \alu_adder_result_ex[22] ;
 wire \alu_adder_result_ex[23] ;
 wire \alu_adder_result_ex[24] ;
 wire \alu_adder_result_ex[25] ;
 wire \alu_adder_result_ex[26] ;
 wire \alu_adder_result_ex[27] ;
 wire \alu_adder_result_ex[28] ;
 wire \alu_adder_result_ex[29] ;
 wire \alu_adder_result_ex[2] ;
 wire \alu_adder_result_ex[30] ;
 wire \alu_adder_result_ex[31] ;
 wire \alu_adder_result_ex[3] ;
 wire \alu_adder_result_ex[4] ;
 wire \alu_adder_result_ex[5] ;
 wire \alu_adder_result_ex[6] ;
 wire \alu_adder_result_ex[7] ;
 wire \alu_adder_result_ex[8] ;
 wire \alu_adder_result_ex[9] ;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net155;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit[0] ;
 wire \cs_registers_i.mcountinhibit[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter[9] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][10] ;
 wire \cs_registers_i.mhpmcounter[2][11] ;
 wire \cs_registers_i.mhpmcounter[2][12] ;
 wire \cs_registers_i.mhpmcounter[2][13] ;
 wire \cs_registers_i.mhpmcounter[2][14] ;
 wire \cs_registers_i.mhpmcounter[2][15] ;
 wire \cs_registers_i.mhpmcounter[2][16] ;
 wire \cs_registers_i.mhpmcounter[2][17] ;
 wire \cs_registers_i.mhpmcounter[2][18] ;
 wire \cs_registers_i.mhpmcounter[2][19] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.mhpmcounter[2][20] ;
 wire \cs_registers_i.mhpmcounter[2][21] ;
 wire \cs_registers_i.mhpmcounter[2][22] ;
 wire \cs_registers_i.mhpmcounter[2][23] ;
 wire \cs_registers_i.mhpmcounter[2][24] ;
 wire \cs_registers_i.mhpmcounter[2][25] ;
 wire \cs_registers_i.mhpmcounter[2][26] ;
 wire \cs_registers_i.mhpmcounter[2][27] ;
 wire \cs_registers_i.mhpmcounter[2][28] ;
 wire \cs_registers_i.mhpmcounter[2][29] ;
 wire \cs_registers_i.mhpmcounter[2][2] ;
 wire \cs_registers_i.mhpmcounter[2][30] ;
 wire \cs_registers_i.mhpmcounter[2][31] ;
 wire \cs_registers_i.mhpmcounter[2][32] ;
 wire \cs_registers_i.mhpmcounter[2][33] ;
 wire \cs_registers_i.mhpmcounter[2][34] ;
 wire \cs_registers_i.mhpmcounter[2][35] ;
 wire \cs_registers_i.mhpmcounter[2][36] ;
 wire \cs_registers_i.mhpmcounter[2][37] ;
 wire \cs_registers_i.mhpmcounter[2][38] ;
 wire \cs_registers_i.mhpmcounter[2][39] ;
 wire \cs_registers_i.mhpmcounter[2][3] ;
 wire \cs_registers_i.mhpmcounter[2][40] ;
 wire \cs_registers_i.mhpmcounter[2][41] ;
 wire \cs_registers_i.mhpmcounter[2][42] ;
 wire \cs_registers_i.mhpmcounter[2][43] ;
 wire \cs_registers_i.mhpmcounter[2][44] ;
 wire \cs_registers_i.mhpmcounter[2][45] ;
 wire \cs_registers_i.mhpmcounter[2][46] ;
 wire \cs_registers_i.mhpmcounter[2][47] ;
 wire \cs_registers_i.mhpmcounter[2][48] ;
 wire \cs_registers_i.mhpmcounter[2][49] ;
 wire \cs_registers_i.mhpmcounter[2][4] ;
 wire \cs_registers_i.mhpmcounter[2][50] ;
 wire \cs_registers_i.mhpmcounter[2][51] ;
 wire \cs_registers_i.mhpmcounter[2][52] ;
 wire \cs_registers_i.mhpmcounter[2][53] ;
 wire \cs_registers_i.mhpmcounter[2][54] ;
 wire \cs_registers_i.mhpmcounter[2][55] ;
 wire \cs_registers_i.mhpmcounter[2][56] ;
 wire \cs_registers_i.mhpmcounter[2][57] ;
 wire \cs_registers_i.mhpmcounter[2][58] ;
 wire \cs_registers_i.mhpmcounter[2][59] ;
 wire \cs_registers_i.mhpmcounter[2][5] ;
 wire \cs_registers_i.mhpmcounter[2][60] ;
 wire \cs_registers_i.mhpmcounter[2][61] ;
 wire \cs_registers_i.mhpmcounter[2][62] ;
 wire \cs_registers_i.mhpmcounter[2][63] ;
 wire \cs_registers_i.mhpmcounter[2][6] ;
 wire \cs_registers_i.mhpmcounter[2][7] ;
 wire \cs_registers_i.mhpmcounter[2][8] ;
 wire \cs_registers_i.mhpmcounter[2][9] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_d[0] ;
 wire \cs_registers_i.mstack_d[1] ;
 wire \cs_registers_i.mstack_d[2] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire \cs_registers_i.priv_lvl_q[1] ;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[24] ;
 wire \load_store_unit_i.rdata_q[25] ;
 wire \load_store_unit_i.rdata_q[26] ;
 wire \load_store_unit_i.rdata_q[27] ;
 wire \load_store_unit_i.rdata_q[28] ;
 wire \load_store_unit_i.rdata_q[29] ;
 wire \load_store_unit_i.rdata_q[30] ;
 wire \load_store_unit_i.rdata_q[31] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net1;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_26_clk_i_regs;
 wire clknet_leaf_27_clk_i_regs;
 wire clknet_leaf_28_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire clknet_leaf_30_clk_i_regs;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_32_clk_i_regs;
 wire clknet_leaf_33_clk_i_regs;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_35_clk_i_regs;
 wire clknet_leaf_36_clk_i_regs;
 wire clknet_leaf_37_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire clknet_leaf_41_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_44_clk_i_regs;
 wire clknet_leaf_45_clk_i_regs;
 wire clknet_leaf_46_clk_i_regs;
 wire clknet_leaf_47_clk_i_regs;
 wire clknet_leaf_48_clk_i_regs;
 wire clknet_leaf_49_clk_i_regs;
 wire clknet_leaf_50_clk_i_regs;
 wire clknet_leaf_51_clk_i_regs;
 wire clknet_leaf_52_clk_i_regs;
 wire clknet_leaf_53_clk_i_regs;
 wire clknet_leaf_54_clk_i_regs;
 wire clknet_leaf_55_clk_i_regs;
 wire clknet_leaf_56_clk_i_regs;
 wire clknet_leaf_57_clk_i_regs;
 wire clknet_leaf_58_clk_i_regs;
 wire clknet_leaf_59_clk_i_regs;
 wire clknet_leaf_60_clk_i_regs;
 wire clknet_leaf_61_clk_i_regs;
 wire clknet_leaf_62_clk_i_regs;
 wire clknet_leaf_63_clk_i_regs;
 wire clknet_leaf_64_clk_i_regs;
 wire clknet_leaf_65_clk_i_regs;
 wire clknet_leaf_66_clk_i_regs;
 wire clknet_leaf_67_clk_i_regs;
 wire clknet_leaf_68_clk_i_regs;
 wire clknet_leaf_69_clk_i_regs;
 wire clknet_leaf_70_clk_i_regs;
 wire clknet_leaf_71_clk_i_regs;
 wire clknet_leaf_72_clk_i_regs;
 wire clknet_leaf_73_clk_i_regs;
 wire clknet_leaf_74_clk_i_regs;
 wire clknet_leaf_75_clk_i_regs;
 wire clknet_leaf_76_clk_i_regs;
 wire clknet_leaf_77_clk_i_regs;
 wire clknet_leaf_78_clk_i_regs;
 wire clknet_leaf_79_clk_i_regs;
 wire clknet_leaf_80_clk_i_regs;
 wire clknet_leaf_81_clk_i_regs;
 wire clknet_leaf_82_clk_i_regs;
 wire clknet_leaf_83_clk_i_regs;
 wire clknet_leaf_84_clk_i_regs;
 wire clknet_leaf_85_clk_i_regs;
 wire clknet_leaf_86_clk_i_regs;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_88_clk_i_regs;
 wire clknet_leaf_89_clk_i_regs;
 wire clknet_leaf_90_clk_i_regs;
 wire clknet_leaf_91_clk_i_regs;
 wire clknet_leaf_92_clk_i_regs;
 wire clknet_leaf_93_clk_i_regs;
 wire clknet_leaf_94_clk_i_regs;
 wire clknet_leaf_95_clk_i_regs;
 wire clknet_leaf_96_clk_i_regs;
 wire clknet_leaf_97_clk_i_regs;
 wire clknet_leaf_98_clk_i_regs;
 wire clknet_leaf_99_clk_i_regs;
 wire clknet_leaf_100_clk_i_regs;
 wire clknet_leaf_101_clk_i_regs;
 wire clknet_leaf_102_clk_i_regs;
 wire clknet_leaf_103_clk_i_regs;
 wire clknet_leaf_104_clk_i_regs;
 wire clknet_leaf_105_clk_i_regs;
 wire clknet_leaf_106_clk_i_regs;
 wire clknet_leaf_107_clk_i_regs;
 wire clknet_leaf_108_clk_i_regs;
 wire clknet_leaf_109_clk_i_regs;
 wire clknet_leaf_110_clk_i_regs;
 wire clknet_leaf_111_clk_i_regs;
 wire clknet_leaf_112_clk_i_regs;
 wire clknet_leaf_113_clk_i_regs;
 wire clknet_leaf_114_clk_i_regs;
 wire clknet_leaf_115_clk_i_regs;
 wire clknet_leaf_116_clk_i_regs;
 wire clknet_leaf_117_clk_i_regs;
 wire clknet_leaf_118_clk_i_regs;
 wire clknet_leaf_119_clk_i_regs;
 wire clknet_leaf_120_clk_i_regs;
 wire clknet_leaf_121_clk_i_regs;
 wire clknet_leaf_122_clk_i_regs;
 wire clknet_leaf_123_clk_i_regs;
 wire clknet_leaf_124_clk_i_regs;
 wire clknet_leaf_125_clk_i_regs;
 wire clknet_leaf_126_clk_i_regs;
 wire clknet_leaf_127_clk_i_regs;
 wire clknet_leaf_128_clk_i_regs;
 wire clknet_leaf_129_clk_i_regs;
 wire clknet_leaf_130_clk_i_regs;
 wire clknet_leaf_131_clk_i_regs;
 wire clknet_leaf_132_clk_i_regs;
 wire clknet_leaf_133_clk_i_regs;
 wire clknet_leaf_134_clk_i_regs;
 wire clknet_leaf_135_clk_i_regs;
 wire clknet_leaf_136_clk_i_regs;
 wire clknet_leaf_137_clk_i_regs;
 wire clknet_leaf_138_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_4_0_0_clk_i_regs;
 wire clknet_4_1_0_clk_i_regs;
 wire clknet_4_2_0_clk_i_regs;
 wire clknet_4_3_0_clk_i_regs;
 wire clknet_4_4_0_clk_i_regs;
 wire clknet_4_5_0_clk_i_regs;
 wire clknet_4_6_0_clk_i_regs;
 wire clknet_4_7_0_clk_i_regs;
 wire clknet_4_8_0_clk_i_regs;
 wire clknet_4_9_0_clk_i_regs;
 wire clknet_4_10_0_clk_i_regs;
 wire clknet_4_11_0_clk_i_regs;
 wire clknet_4_12_0_clk_i_regs;
 wire clknet_4_13_0_clk_i_regs;
 wire clknet_4_14_0_clk_i_regs;
 wire clknet_4_15_0_clk_i_regs;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net392;
 wire net393;
 wire net397;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net440;
 wire net441;
 wire net442;
 wire net444;
 wire net445;
 wire net447;
 wire net448;
 wire net449;
 wire net450;

 BUF_X4 _16113_ (.A(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_10287_));
 INV_X2 _16114_ (.A(_10287_),
    .ZN(_10288_));
 BUF_X8 _16115_ (.A(_10288_),
    .Z(_10289_));
 BUF_X2 _16116_ (.A(\id_stage_i.controller_i.instr_i[1] ),
    .Z(_10290_));
 BUF_X2 _16117_ (.A(\id_stage_i.controller_i.instr_i[0] ),
    .Z(_10291_));
 NAND2_X4 _16118_ (.A1(_10290_),
    .A2(_10291_),
    .ZN(_10292_));
 BUF_X8 _16119_ (.A(\id_stage_i.controller_i.instr_i[3] ),
    .Z(_10293_));
 BUF_X1 rebuffer28 (.A(_10323_),
    .Z(net299));
 OR2_X4 _16121_ (.A1(_10293_),
    .A2(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_10295_));
 BUF_X8 _16122_ (.A(_10295_),
    .Z(_10296_));
 NOR3_X2 _16123_ (.A1(_10289_),
    .A2(_10292_),
    .A3(_10296_),
    .ZN(_10297_));
 BUF_X2 _16124_ (.A(\id_stage_i.controller_i.instr_i[6] ),
    .Z(_10298_));
 BUF_X4 _16125_ (.A(_10298_),
    .Z(_10299_));
 BUF_X8 _16126_ (.A(\id_stage_i.controller_i.instr_i[4] ),
    .Z(_10300_));
 BUF_X2 _16127_ (.A(_00172_),
    .Z(_10301_));
 NOR2_X4 _16128_ (.A1(_10300_),
    .A2(_10301_),
    .ZN(_10302_));
 NOR2_X1 _16129_ (.A1(_10299_),
    .A2(_10302_),
    .ZN(_10303_));
 BUF_X4 _16130_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .Z(_10304_));
 INV_X4 _16131_ (.A(_10304_),
    .ZN(_10305_));
 BUF_X4 _16132_ (.A(\id_stage_i.id_fsm_q ),
    .Z(_10306_));
 OR2_X4 _16133_ (.A1(net310),
    .A2(_10301_),
    .ZN(_10307_));
 NOR3_X2 _16134_ (.A1(_10305_),
    .A2(_10306_),
    .A3(_10307_),
    .ZN(_10308_));
 BUF_X8 _16135_ (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_10309_));
 BUF_X16 _16136_ (.A(_10309_),
    .Z(_10310_));
 AND2_X1 _16137_ (.A1(_10290_),
    .A2(_10291_),
    .ZN(_10311_));
 BUF_X4 _16138_ (.A(_10311_),
    .Z(_10312_));
 NOR2_X4 _16139_ (.A1(_10293_),
    .A2(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_10313_));
 NOR2_X4 _16140_ (.A1(_10300_),
    .A2(_10299_),
    .ZN(_10314_));
 NAND3_X4 _16141_ (.A1(_10312_),
    .A2(_10313_),
    .A3(_10314_),
    .ZN(_10315_));
 OAI221_X2 _16142_ (.A(_10297_),
    .B1(_10303_),
    .B2(_10308_),
    .C1(_10310_),
    .C2(_10315_),
    .ZN(_10316_));
 BUF_X8 _16143_ (.A(_10316_),
    .Z(_10317_));
 INV_X1 _16144_ (.A(_16085_),
    .ZN(_10318_));
 BUF_X4 _16145_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .Z(_10319_));
 BUF_X2 _16146_ (.A(_00171_),
    .Z(_10320_));
 AND2_X1 _16147_ (.A1(_10319_),
    .A2(_10320_),
    .ZN(_10321_));
 BUF_X1 _16148_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .Z(_10322_));
 MUX2_X1 _16149_ (.A(_10322_),
    .B(_10320_),
    .S(_10319_),
    .Z(_10323_));
 CLKBUF_X3 _16150_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .Z(_10324_));
 INV_X2 _16151_ (.A(_10324_),
    .ZN(_10325_));
 AOI22_X4 _16152_ (.A1(_10318_),
    .A2(_10321_),
    .B1(net299),
    .B2(_10325_),
    .ZN(_10326_));
 INV_X2 _16153_ (.A(_10293_),
    .ZN(_10327_));
 INV_X2 _16154_ (.A(_10298_),
    .ZN(_10328_));
 AND3_X1 _16155_ (.A1(_10290_),
    .A2(_10291_),
    .A3(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_10329_));
 BUF_X4 _16156_ (.A(_10329_),
    .Z(_10330_));
 NAND4_X4 _16157_ (.A1(_10327_),
    .A2(net311),
    .A3(_10328_),
    .A4(_10330_),
    .ZN(_10331_));
 NAND4_X4 _16158_ (.A1(_10312_),
    .A2(_10287_),
    .A3(_10313_),
    .A4(_10302_),
    .ZN(_10332_));
 NOR2_X4 _16159_ (.A1(_10305_),
    .A2(_10306_),
    .ZN(_10333_));
 OAI211_X4 _16160_ (.A(_10326_),
    .B(_10331_),
    .C1(_10332_),
    .C2(_10333_),
    .ZN(_10334_));
 BUF_X8 _16161_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(_10335_));
 INV_X2 _16162_ (.A(_10335_),
    .ZN(_10336_));
 BUF_X4 _16163_ (.A(_10336_),
    .Z(_10337_));
 BUF_X4 _16164_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_10338_));
 NAND3_X2 _16165_ (.A1(_10290_),
    .A2(_10291_),
    .A3(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_10339_));
 BUF_X4 _16166_ (.A(_10339_),
    .Z(_10340_));
 BUF_X4 _16167_ (.A(_10293_),
    .Z(_10341_));
 AND3_X2 _16168_ (.A1(_10341_),
    .A2(_10289_),
    .A3(_10314_),
    .ZN(_10342_));
 BUF_X2 _16169_ (.A(\id_stage_i.controller_i.instr_i[13] ),
    .Z(_10343_));
 BUF_X4 _16170_ (.A(_10343_),
    .Z(_10344_));
 BUF_X2 _16171_ (.A(\id_stage_i.controller_i.instr_i[12] ),
    .Z(_10345_));
 INV_X4 _16172_ (.A(_10345_),
    .ZN(_10346_));
 BUF_X4 _16173_ (.A(_00173_),
    .Z(_10347_));
 INV_X4 _16174_ (.A(_10347_),
    .ZN(_10348_));
 NOR3_X4 _16175_ (.A1(_10344_),
    .A2(_10346_),
    .A3(_10348_),
    .ZN(_10349_));
 INV_X4 _16176_ (.A(_10306_),
    .ZN(_10350_));
 NAND3_X1 _16177_ (.A1(_10327_),
    .A2(_10304_),
    .A3(_10350_),
    .ZN(_10351_));
 NOR2_X4 _16178_ (.A1(_10289_),
    .A2(_10307_),
    .ZN(_10352_));
 AOI22_X2 _16179_ (.A1(_10342_),
    .A2(_10349_),
    .B1(_10351_),
    .B2(_10352_),
    .ZN(_10353_));
 NOR2_X1 _16180_ (.A1(_10340_),
    .A2(_10353_),
    .ZN(_10354_));
 NAND2_X1 _16181_ (.A1(_10338_),
    .A2(_10354_),
    .ZN(_10355_));
 AND2_X1 _16182_ (.A1(_10325_),
    .A2(_10323_),
    .ZN(_10356_));
 NAND2_X1 _16183_ (.A1(_10319_),
    .A2(_10320_),
    .ZN(_10357_));
 NOR2_X1 _16184_ (.A1(_16085_),
    .A2(_10357_),
    .ZN(_10358_));
 OR2_X1 _16185_ (.A1(_10356_),
    .A2(_10358_),
    .ZN(_10359_));
 BUF_X4 _16186_ (.A(_10359_),
    .Z(_10360_));
 BUF_X4 _16187_ (.A(_10360_),
    .Z(_10361_));
 MUX2_X1 _16188_ (.A(_10298_),
    .B(_10301_),
    .S(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_10362_));
 NOR3_X2 _16189_ (.A1(net311),
    .A2(_10340_),
    .A3(_10362_),
    .ZN(_10363_));
 INV_X1 _16190_ (.A(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_10364_));
 NOR2_X1 _16191_ (.A1(_10327_),
    .A2(_10364_),
    .ZN(_10365_));
 NOR3_X2 _16192_ (.A1(_10341_),
    .A2(_10289_),
    .A3(_10301_),
    .ZN(_10366_));
 OAI211_X2 _16193_ (.A(_10312_),
    .B(_10363_),
    .C1(_10365_),
    .C2(_10366_),
    .ZN(_10367_));
 NAND2_X4 _16194_ (.A1(_10304_),
    .A2(_10350_),
    .ZN(_10368_));
 AOI22_X2 _16195_ (.A1(_10368_),
    .A2(_10352_),
    .B1(_10342_),
    .B2(_10349_),
    .ZN(_10369_));
 OR3_X1 _16196_ (.A1(_10360_),
    .A2(_10367_),
    .A3(_10369_),
    .ZN(_10370_));
 BUF_X4 _16197_ (.A(_10370_),
    .Z(_10371_));
 INV_X2 _16198_ (.A(_10300_),
    .ZN(_10372_));
 NOR4_X4 _16199_ (.A1(_10339_),
    .A2(_10372_),
    .A3(_10298_),
    .A4(_10293_),
    .ZN(_10373_));
 NOR3_X4 _16200_ (.A1(_10289_),
    .A2(_10310_),
    .A3(_10315_),
    .ZN(_10374_));
 NOR2_X4 _16201_ (.A1(_10373_),
    .A2(_10374_),
    .ZN(_10375_));
 AOI21_X1 _16202_ (.A(_10361_),
    .B1(_10371_),
    .B2(_10375_),
    .ZN(_10376_));
 MUX2_X1 _16203_ (.A(_10337_),
    .B(_10355_),
    .S(_10376_),
    .Z(_10377_));
 NAND3_X2 _16204_ (.A1(_10293_),
    .A2(_10288_),
    .A3(_10314_),
    .ZN(_10378_));
 INV_X1 _16205_ (.A(_10344_),
    .ZN(_10379_));
 BUF_X4 _16206_ (.A(_10379_),
    .Z(_10380_));
 BUF_X4 _16207_ (.A(_10345_),
    .Z(_10381_));
 NAND3_X2 _16208_ (.A1(_10380_),
    .A2(_10381_),
    .A3(_10347_),
    .ZN(_10382_));
 NOR3_X2 _16209_ (.A1(_10341_),
    .A2(_10305_),
    .A3(_10306_),
    .ZN(_10383_));
 NAND2_X2 _16210_ (.A1(_10287_),
    .A2(_10302_),
    .ZN(_10384_));
 OAI22_X4 _16211_ (.A1(_10378_),
    .A2(_10382_),
    .B1(_10383_),
    .B2(_10384_),
    .ZN(_10385_));
 AOI21_X4 _16212_ (.A(_10360_),
    .B1(_10330_),
    .B2(_10385_),
    .ZN(_10386_));
 AOI21_X4 _16213_ (.A(_10334_),
    .B1(_10371_),
    .B2(_10375_),
    .ZN(_10387_));
 OAI21_X2 _16214_ (.A(_10331_),
    .B1(_10332_),
    .B2(_10333_),
    .ZN(_10388_));
 NOR2_X4 _16215_ (.A1(_10360_),
    .A2(_10388_),
    .ZN(_10389_));
 NAND2_X1 _16216_ (.A1(net311),
    .A2(_10328_),
    .ZN(_10390_));
 OAI33_X1 _16217_ (.A1(_10341_),
    .A2(_10390_),
    .A3(_10340_),
    .B1(_10360_),
    .B2(_10369_),
    .B3(_10367_),
    .ZN(_10391_));
 NOR3_X4 _16218_ (.A1(_10389_),
    .A2(_10374_),
    .A3(net20),
    .ZN(_10392_));
 OAI21_X2 _16219_ (.A(_10386_),
    .B1(_10387_),
    .B2(_10392_),
    .ZN(_10393_));
 BUF_X4 _16220_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .Z(_10394_));
 INV_X1 _16221_ (.A(_10394_),
    .ZN(_10395_));
 OAI221_X2 _16222_ (.A(_10317_),
    .B1(_10334_),
    .B2(_10377_),
    .C1(_10393_),
    .C2(_10395_),
    .ZN(_10396_));
 BUF_X4 _16223_ (.A(_10361_),
    .Z(_10397_));
 BUF_X4 _16224_ (.A(_10397_),
    .Z(_10398_));
 OAI21_X2 _16225_ (.A(_10297_),
    .B1(_10303_),
    .B2(_10308_),
    .ZN(_10399_));
 NOR2_X1 _16226_ (.A1(_10292_),
    .A2(_10296_),
    .ZN(_10400_));
 AND2_X2 _16227_ (.A1(_10400_),
    .A2(_10314_),
    .ZN(_10401_));
 INV_X4 _16228_ (.A(_10309_),
    .ZN(_10402_));
 AOI21_X4 _16229_ (.A(_10399_),
    .B1(_10401_),
    .B2(_10402_),
    .ZN(_10403_));
 BUF_X4 _16230_ (.A(_10335_),
    .Z(_10404_));
 BUF_X8 _16231_ (.A(_10404_),
    .Z(_10405_));
 BUF_X8 _16232_ (.A(_10405_),
    .Z(_10406_));
 MUX2_X1 _16233_ (.A(_00163_),
    .B(_00165_),
    .S(_10406_),
    .Z(_10407_));
 BUF_X8 _16234_ (.A(_10335_),
    .Z(_10408_));
 BUF_X8 _16235_ (.A(_10408_),
    .Z(_10409_));
 BUF_X4 _16236_ (.A(_10409_),
    .Z(_10410_));
 MUX2_X1 _16237_ (.A(_00164_),
    .B(_00166_),
    .S(_10410_),
    .Z(_10411_));
 BUF_X8 _16238_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(_10412_));
 BUF_X8 _16239_ (.A(_10412_),
    .Z(_10413_));
 BUF_X4 _16240_ (.A(_10413_),
    .Z(_10414_));
 MUX2_X1 _16241_ (.A(_10407_),
    .B(_10411_),
    .S(_10414_),
    .Z(_10415_));
 MUX2_X1 _16242_ (.A(_00155_),
    .B(_00157_),
    .S(_10410_),
    .Z(_10416_));
 MUX2_X1 _16243_ (.A(_00156_),
    .B(_00158_),
    .S(_10410_),
    .Z(_10417_));
 MUX2_X1 _16244_ (.A(_10416_),
    .B(_10417_),
    .S(_10414_),
    .Z(_10418_));
 BUF_X4 _16245_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(_10419_));
 INV_X2 _16246_ (.A(_10419_),
    .ZN(_10420_));
 BUF_X8 _16247_ (.A(_10420_),
    .Z(_10421_));
 MUX2_X1 _16248_ (.A(_10415_),
    .B(_10418_),
    .S(_10421_),
    .Z(_10422_));
 MUX2_X1 _16249_ (.A(_00167_),
    .B(_00169_),
    .S(_10410_),
    .Z(_10423_));
 MUX2_X1 _16250_ (.A(_00168_),
    .B(_00170_),
    .S(_10410_),
    .Z(_10424_));
 MUX2_X1 _16251_ (.A(_10423_),
    .B(_10424_),
    .S(_10414_),
    .Z(_10425_));
 MUX2_X1 _16252_ (.A(_00159_),
    .B(_00161_),
    .S(_10410_),
    .Z(_10426_));
 MUX2_X1 _16253_ (.A(_00160_),
    .B(_00162_),
    .S(_10410_),
    .Z(_10427_));
 MUX2_X1 _16254_ (.A(_10426_),
    .B(_10427_),
    .S(_10414_),
    .Z(_10428_));
 MUX2_X1 _16255_ (.A(_10425_),
    .B(_10428_),
    .S(_10421_),
    .Z(_10429_));
 BUF_X4 _16256_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(_10430_));
 BUF_X4 _16257_ (.A(_10430_),
    .Z(_10431_));
 BUF_X8 _16258_ (.A(_10431_),
    .Z(_10432_));
 MUX2_X1 _16259_ (.A(_10422_),
    .B(_10429_),
    .S(_10432_),
    .Z(_10433_));
 BUF_X4 _16260_ (.A(_10430_),
    .Z(_10434_));
 INV_X4 _16261_ (.A(_10434_),
    .ZN(_10435_));
 BUF_X4 _16262_ (.A(_10435_),
    .Z(_10436_));
 BUF_X4 _16263_ (.A(_10404_),
    .Z(_10437_));
 BUF_X8 _16264_ (.A(_10437_),
    .Z(_10438_));
 BUF_X8 _16265_ (.A(_10438_),
    .Z(_10439_));
 MUX2_X1 _16266_ (.A(_00151_),
    .B(_00153_),
    .S(_10439_),
    .Z(_10440_));
 MUX2_X1 _16267_ (.A(_00152_),
    .B(_00154_),
    .S(_10439_),
    .Z(_10441_));
 BUF_X4 _16268_ (.A(_10412_),
    .Z(_10442_));
 BUF_X4 _16269_ (.A(_10442_),
    .Z(_10443_));
 BUF_X4 _16270_ (.A(_10443_),
    .Z(_10444_));
 MUX2_X1 _16271_ (.A(_10440_),
    .B(_10441_),
    .S(_10444_),
    .Z(_10445_));
 MUX2_X1 _16272_ (.A(_00143_),
    .B(_00145_),
    .S(_10439_),
    .Z(_10446_));
 MUX2_X1 _16273_ (.A(_00144_),
    .B(_00146_),
    .S(_10439_),
    .Z(_10447_));
 MUX2_X1 _16274_ (.A(_10446_),
    .B(_10447_),
    .S(_10444_),
    .Z(_10448_));
 MUX2_X1 _16275_ (.A(_10445_),
    .B(_10448_),
    .S(_10421_),
    .Z(_10449_));
 NOR2_X1 _16276_ (.A1(_10436_),
    .A2(_10449_),
    .ZN(_10450_));
 BUF_X8 _16277_ (.A(_10419_),
    .Z(_10451_));
 BUF_X4 _16278_ (.A(_10408_),
    .Z(_10452_));
 BUF_X4 _16279_ (.A(_10452_),
    .Z(_10453_));
 BUF_X4 _16280_ (.A(_10453_),
    .Z(_10454_));
 NOR2_X1 _16281_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A2(_10454_),
    .ZN(_10455_));
 BUF_X32 _16282_ (.A(net432),
    .Z(_10456_));
 BUF_X32 _16283_ (.A(_10456_),
    .Z(_10457_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 BUF_X32 _16285_ (.A(_10457_),
    .Z(_10459_));
 AOI21_X1 _16286_ (.A(_10455_),
    .B1(net357),
    .B2(_00142_),
    .ZN(_10460_));
 NOR2_X1 _16287_ (.A1(_10444_),
    .A2(_00141_),
    .ZN(_10461_));
 AOI221_X2 _16288_ (.A(_10451_),
    .B1(_10460_),
    .B2(_10444_),
    .C1(_10461_),
    .C2(net357),
    .ZN(_10462_));
 MUX2_X1 _16289_ (.A(_00147_),
    .B(_00149_),
    .S(net357),
    .Z(_10463_));
 MUX2_X1 _16290_ (.A(_00148_),
    .B(_00150_),
    .S(net357),
    .Z(_10464_));
 BUF_X8 _16291_ (.A(_10413_),
    .Z(_10465_));
 BUF_X8 _16292_ (.A(_10465_),
    .Z(_10466_));
 MUX2_X1 _16293_ (.A(_10463_),
    .B(_10464_),
    .S(_10466_),
    .Z(_10467_));
 BUF_X8 _16294_ (.A(_10451_),
    .Z(_10468_));
 AOI21_X1 _16295_ (.A(_10462_),
    .B1(_10467_),
    .B2(_10468_),
    .ZN(_10469_));
 AOI21_X2 _16296_ (.A(_10450_),
    .B1(_10469_),
    .B2(_10436_),
    .ZN(_10470_));
 BUF_X4 _16297_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(_10471_));
 INV_X8 _16298_ (.A(_10471_),
    .ZN(_10472_));
 BUF_X4 _16299_ (.A(_10472_),
    .Z(_10473_));
 BUF_X8 _16300_ (.A(_10473_),
    .Z(_10474_));
 MUX2_X2 _16301_ (.A(_10433_),
    .B(_10470_),
    .S(_10474_),
    .Z(_10475_));
 AOI21_X4 _16302_ (.A(_10398_),
    .B1(_10403_),
    .B2(_10475_),
    .ZN(_10476_));
 NAND2_X4 _16303_ (.A1(_10396_),
    .A2(_10476_),
    .ZN(_15834_));
 INV_X2 _16304_ (.A(_15834_),
    .ZN(_15846_));
 CLKBUF_X3 _16305_ (.A(_10381_),
    .Z(_10477_));
 NOR2_X1 _16306_ (.A1(_10477_),
    .A2(_10348_),
    .ZN(_10478_));
 NOR2_X4 _16307_ (.A1(_10368_),
    .A2(_10332_),
    .ZN(_10479_));
 NAND2_X4 _16308_ (.A1(_10312_),
    .A2(_10313_),
    .ZN(_10480_));
 NAND3_X4 _16309_ (.A1(_10300_),
    .A2(_10288_),
    .A3(_10328_),
    .ZN(_10481_));
 NAND2_X2 _16310_ (.A1(_10309_),
    .A2(_10345_),
    .ZN(_10482_));
 NAND2_X1 _16311_ (.A1(_10343_),
    .A2(_10347_),
    .ZN(_10483_));
 NOR2_X2 _16312_ (.A1(_10482_),
    .A2(_10483_),
    .ZN(_10484_));
 INV_X1 _16313_ (.A(_00176_),
    .ZN(_10485_));
 AOI211_X2 _16314_ (.A(_10343_),
    .B(_10485_),
    .C1(_10346_),
    .C2(_10309_),
    .ZN(_10486_));
 NOR4_X4 _16315_ (.A1(_10480_),
    .A2(_10481_),
    .A3(_10484_),
    .A4(_10486_),
    .ZN(_10487_));
 BUF_X4 _16316_ (.A(_10344_),
    .Z(_10488_));
 MUX2_X1 _16317_ (.A(_10479_),
    .B(_10487_),
    .S(_10488_),
    .Z(_10489_));
 NAND2_X2 _16318_ (.A1(_10344_),
    .A2(_10346_),
    .ZN(_10490_));
 OAI33_X1 _16319_ (.A1(_10488_),
    .A2(_10368_),
    .A3(_10332_),
    .B1(_10481_),
    .B2(_10490_),
    .B3(_10480_),
    .ZN(_10491_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 BUF_X16 _16321_ (.A(_10310_),
    .Z(_10493_));
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 BUF_X8 _16323_ (.A(_10493_),
    .Z(_10495_));
 AOI22_X1 _16324_ (.A1(_10478_),
    .A2(_10489_),
    .B1(_10491_),
    .B2(_10495_),
    .ZN(_10496_));
 BUF_X2 _16325_ (.A(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_10497_));
 BUF_X4 _16326_ (.A(_10497_),
    .Z(_10498_));
 INV_X1 _16327_ (.A(_10498_),
    .ZN(_10499_));
 BUF_X4 _16328_ (.A(\id_stage_i.controller_i.instr_i[27] ),
    .Z(_10500_));
 BUF_X8 _16329_ (.A(\id_stage_i.controller_i.instr_i[28] ),
    .Z(_10501_));
 BUF_X4 _16330_ (.A(\id_stage_i.controller_i.instr_i[29] ),
    .Z(_10502_));
 INV_X1 _16331_ (.A(_00174_),
    .ZN(_10503_));
 NOR4_X2 _16332_ (.A1(_10500_),
    .A2(_10501_),
    .A3(_10502_),
    .A4(_10503_),
    .ZN(_10504_));
 AND4_X1 _16333_ (.A1(_10310_),
    .A2(_10380_),
    .A3(_10381_),
    .A4(_10504_),
    .ZN(_10505_));
 NAND3_X1 _16334_ (.A1(_10499_),
    .A2(_10487_),
    .A3(_10505_),
    .ZN(_10506_));
 BUF_X2 _16335_ (.A(\id_stage_i.controller_i.instr_i[25] ),
    .Z(_10507_));
 INV_X4 _16336_ (.A(_10507_),
    .ZN(_10508_));
 BUF_X4 _16337_ (.A(\id_stage_i.controller_i.instr_i[31] ),
    .Z(_10509_));
 INV_X2 _16338_ (.A(_10509_),
    .ZN(_10510_));
 NOR4_X4 _16339_ (.A1(_10500_),
    .A2(_10502_),
    .A3(_10501_),
    .A4(\id_stage_i.controller_i.instr_i[26] ),
    .ZN(_10511_));
 NAND3_X2 _16340_ (.A1(_10508_),
    .A2(_10510_),
    .A3(net282),
    .ZN(_10512_));
 NAND2_X2 _16341_ (.A1(_10300_),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .ZN(_10513_));
 NOR4_X4 _16342_ (.A1(_10296_),
    .A2(_10292_),
    .A3(_10299_),
    .A4(_10513_),
    .ZN(_10514_));
 NOR2_X1 _16343_ (.A1(_10498_),
    .A2(_10482_),
    .ZN(_10515_));
 NOR3_X2 _16344_ (.A1(_10495_),
    .A2(_10381_),
    .A3(_10499_),
    .ZN(_10516_));
 OAI21_X1 _16345_ (.A(_10380_),
    .B1(_10515_),
    .B2(_10516_),
    .ZN(_10517_));
 OAI21_X1 _16346_ (.A(_10517_),
    .B1(_10490_),
    .B2(_10498_),
    .ZN(_10518_));
 NAND2_X1 _16347_ (.A1(_10514_),
    .A2(_10518_),
    .ZN(_10519_));
 OR2_X2 _16348_ (.A1(_10512_),
    .A2(_10519_),
    .ZN(_10520_));
 AND3_X4 _16349_ (.A1(_10496_),
    .A2(_10506_),
    .A3(_10520_),
    .ZN(_15357_));
 INV_X4 _16350_ (.A(_15357_),
    .ZN(_15364_));
 AOI21_X1 _16351_ (.A(_10488_),
    .B1(_10348_),
    .B2(_10504_),
    .ZN(_10521_));
 BUF_X4 _16352_ (.A(_10347_),
    .Z(_10522_));
 OAI21_X1 _16353_ (.A(_10477_),
    .B1(_10522_),
    .B2(_10488_),
    .ZN(_10523_));
 INV_X1 _16354_ (.A(_10523_),
    .ZN(_10524_));
 OAI221_X2 _16355_ (.A(_10487_),
    .B1(_10521_),
    .B2(_10482_),
    .C1(_10524_),
    .C2(_10495_),
    .ZN(_10525_));
 NOR2_X2 _16356_ (.A1(_10488_),
    .A2(_10346_),
    .ZN(_10526_));
 INV_X1 _16357_ (.A(_10490_),
    .ZN(_10527_));
 OAI21_X1 _16358_ (.A(_10495_),
    .B1(_10526_),
    .B2(_10527_),
    .ZN(_10528_));
 NAND3_X1 _16359_ (.A1(_10382_),
    .A2(_10479_),
    .A3(_10528_),
    .ZN(_10529_));
 NOR4_X4 _16360_ (.A1(_10327_),
    .A2(net311),
    .A3(_10340_),
    .A4(_10362_),
    .ZN(_10530_));
 NOR3_X2 _16361_ (.A1(_10299_),
    .A2(_10292_),
    .A3(_10296_),
    .ZN(_10531_));
 NOR4_X4 _16362_ (.A1(_10293_),
    .A2(_10288_),
    .A3(_10292_),
    .A4(_10307_),
    .ZN(_10532_));
 NOR4_X4 _16363_ (.A1(_10373_),
    .A2(_10530_),
    .A3(_10531_),
    .A4(_10532_),
    .ZN(_10533_));
 NOR2_X2 _16364_ (.A1(_10287_),
    .A2(_10299_),
    .ZN(_10534_));
 AND4_X2 _16365_ (.A1(_10341_),
    .A2(_10372_),
    .A3(_10330_),
    .A4(_10534_),
    .ZN(_10535_));
 NAND2_X2 _16366_ (.A1(_10380_),
    .A2(_10522_),
    .ZN(_10536_));
 AOI21_X2 _16367_ (.A(_10533_),
    .B1(_10535_),
    .B2(_10536_),
    .ZN(_10537_));
 CLKBUF_X2 _16368_ (.A(_00177_),
    .Z(_10538_));
 INV_X1 _16369_ (.A(_10538_),
    .ZN(_10539_));
 NOR2_X2 _16370_ (.A1(_10509_),
    .A2(_10497_),
    .ZN(_10540_));
 NAND2_X2 _16371_ (.A1(_10511_),
    .A2(_10540_),
    .ZN(_10541_));
 AOI21_X1 _16372_ (.A(_10507_),
    .B1(_10346_),
    .B2(net315),
    .ZN(_10542_));
 AOI211_X2 _16373_ (.A(_10507_),
    .B(_10509_),
    .C1(_10497_),
    .C2(_10343_),
    .ZN(_10543_));
 NAND2_X1 _16374_ (.A1(_10543_),
    .A2(_10511_),
    .ZN(_10544_));
 NOR2_X1 _16375_ (.A1(_10344_),
    .A2(_10497_),
    .ZN(_10545_));
 NOR3_X1 _16376_ (.A1(_10309_),
    .A2(_10346_),
    .A3(_10545_),
    .ZN(_10546_));
 OAI21_X1 _16377_ (.A(_10538_),
    .B1(_10381_),
    .B2(_10402_),
    .ZN(_10547_));
 OAI33_X1 _16378_ (.A1(_10541_),
    .A2(_10539_),
    .A3(_10542_),
    .B1(_10544_),
    .B2(_10546_),
    .B3(_10547_),
    .ZN(_10548_));
 NAND2_X2 _16379_ (.A1(_10379_),
    .A2(_10381_),
    .ZN(_10549_));
 MUX2_X1 _16380_ (.A(_10381_),
    .B(_10549_),
    .S(_10402_),
    .Z(_10550_));
 NAND3_X1 _16381_ (.A1(_10508_),
    .A2(_10511_),
    .A3(_10540_),
    .ZN(_10551_));
 OAI21_X4 _16382_ (.A(net277),
    .B1(_10550_),
    .B2(_10551_),
    .ZN(_10552_));
 NAND2_X4 _16383_ (.A1(_10514_),
    .A2(_10552_),
    .ZN(_10553_));
 NAND4_X4 _16384_ (.A1(_10525_),
    .A2(_10553_),
    .A3(_10537_),
    .A4(_10529_),
    .ZN(_15358_));
 INV_X4 _16385_ (.A(_15358_),
    .ZN(_15361_));
 NOR2_X1 _16386_ (.A1(_10344_),
    .A2(_10348_),
    .ZN(_10554_));
 NAND4_X4 _16387_ (.A1(_10341_),
    .A2(_10372_),
    .A3(_10330_),
    .A4(_10534_),
    .ZN(_10555_));
 NAND3_X2 _16388_ (.A1(net311),
    .A2(_10287_),
    .A3(_10299_),
    .ZN(_10556_));
 OR3_X4 _16389_ (.A1(_10292_),
    .A2(_10296_),
    .A3(_10556_),
    .ZN(_10557_));
 OAI221_X2 _16390_ (.A(_10326_),
    .B1(_10554_),
    .B2(_10555_),
    .C1(_10557_),
    .C2(_10522_),
    .ZN(_10558_));
 NOR4_X1 _16391_ (.A1(_10327_),
    .A2(_10289_),
    .A3(_10307_),
    .A4(_10340_),
    .ZN(_10559_));
 AOI21_X2 _16392_ (.A(_10559_),
    .B1(_10373_),
    .B2(_10289_),
    .ZN(_10560_));
 NAND2_X1 _16393_ (.A1(_10299_),
    .A2(_10513_),
    .ZN(_10561_));
 AOI221_X2 _16394_ (.A(_10532_),
    .B1(_10561_),
    .B2(_10400_),
    .C1(_10330_),
    .C2(_10342_),
    .ZN(_10562_));
 AOI21_X4 _16395_ (.A(_10558_),
    .B1(_10560_),
    .B2(_10562_),
    .ZN(_10563_));
 BUF_X2 _16396_ (.A(_10563_),
    .Z(_10564_));
 BUF_X4 _16397_ (.A(_10564_),
    .Z(_10565_));
 BUF_X4 _16398_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .Z(_10566_));
 INV_X8 _16399_ (.A(_10566_),
    .ZN(_10567_));
 BUF_X4 _16400_ (.A(_10567_),
    .Z(_10568_));
 BUF_X4 _16401_ (.A(_10568_),
    .Z(_10569_));
 BUF_X4 _16402_ (.A(_10569_),
    .Z(_10570_));
 BUF_X4 _16403_ (.A(_10570_),
    .Z(_10571_));
 BUF_X4 _16404_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .Z(_10572_));
 INV_X4 _16405_ (.A(_10572_),
    .ZN(_10573_));
 BUF_X8 _16406_ (.A(_10573_),
    .Z(_10574_));
 BUF_X4 _16407_ (.A(_10574_),
    .Z(_10575_));
 BUF_X4 _16408_ (.A(_10575_),
    .Z(_10576_));
 BUF_X4 _16409_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(_10577_));
 INV_X1 _16410_ (.A(_10577_),
    .ZN(_10578_));
 BUF_X4 _16411_ (.A(_10578_),
    .Z(_10579_));
 BUF_X8 _16412_ (.A(_10579_),
    .Z(_10580_));
 BUF_X4 _16413_ (.A(_10580_),
    .Z(_10581_));
 BUF_X4 _16414_ (.A(_10581_),
    .Z(_10582_));
 BUF_X4 _16415_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(_10583_));
 BUF_X8 _16416_ (.A(_10583_),
    .Z(_10584_));
 BUF_X8 _16417_ (.A(_10584_),
    .Z(_10585_));
 BUF_X4 rebuffer87 (.A(_12683_),
    .Z(net358));
 BUF_X8 _16419_ (.A(_10585_),
    .Z(_10587_));
 BUF_X4 _16420_ (.A(_10587_),
    .Z(_10588_));
 BUF_X4 _16421_ (.A(_10588_),
    .Z(_10589_));
 MUX2_X1 _16422_ (.A(_00156_),
    .B(_00158_),
    .S(_10589_),
    .Z(_10590_));
 NOR2_X1 _16423_ (.A1(_10582_),
    .A2(_10590_),
    .ZN(_10591_));
 BUF_X8 _16424_ (.A(_10577_),
    .Z(_10592_));
 BUF_X8 _16425_ (.A(_10592_),
    .Z(_10593_));
 BUF_X8 _16426_ (.A(_10593_),
    .Z(_10594_));
 BUF_X8 _16427_ (.A(_10594_),
    .Z(_10595_));
 BUF_X4 _16428_ (.A(_10595_),
    .Z(_10596_));
 BUF_X4 _16429_ (.A(_10596_),
    .Z(_10597_));
 BUF_X8 _16430_ (.A(_10584_),
    .Z(_10598_));
 BUF_X8 _16431_ (.A(_10598_),
    .Z(_10599_));
 BUF_X8 _16432_ (.A(_10599_),
    .Z(_10600_));
 BUF_X4 _16433_ (.A(_10600_),
    .Z(_10601_));
 BUF_X8 _16434_ (.A(_10601_),
    .Z(_10602_));
 MUX2_X1 _16435_ (.A(_00155_),
    .B(_00157_),
    .S(_10602_),
    .Z(_10603_));
 NOR2_X1 _16436_ (.A1(_10597_),
    .A2(_10603_),
    .ZN(_10604_));
 NOR3_X2 _16437_ (.A1(_10576_),
    .A2(_10591_),
    .A3(_10604_),
    .ZN(_10605_));
 BUF_X8 _16438_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(_10606_));
 INV_X4 _16439_ (.A(_10606_),
    .ZN(_10607_));
 BUF_X8 _16440_ (.A(_10607_),
    .Z(_10608_));
 BUF_X8 _16441_ (.A(_10608_),
    .Z(_10609_));
 BUF_X4 _16442_ (.A(_10609_),
    .Z(_10610_));
 BUF_X4 _16443_ (.A(_10583_),
    .Z(_10611_));
 BUF_X4 _16444_ (.A(_10611_),
    .Z(_10612_));
 BUF_X4 _16445_ (.A(_10612_),
    .Z(_10613_));
 BUF_X4 _16446_ (.A(_10613_),
    .Z(_10614_));
 BUF_X4 _16447_ (.A(_10614_),
    .Z(_10615_));
 BUF_X4 _16448_ (.A(_10615_),
    .Z(_10616_));
 NOR2_X1 _16449_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A2(_10616_),
    .ZN(_10617_));
 BUF_X4 _16450_ (.A(_10584_),
    .Z(_10618_));
 BUF_X4 _16451_ (.A(_10618_),
    .Z(_10619_));
 BUF_X4 _16452_ (.A(_10619_),
    .Z(_10620_));
 BUF_X8 _16453_ (.A(_10620_),
    .Z(_10621_));
 BUF_X8 _16454_ (.A(_10621_),
    .Z(_10622_));
 AND2_X1 _16455_ (.A1(_00142_),
    .A2(_10622_),
    .ZN(_10623_));
 NOR3_X1 _16456_ (.A1(_10582_),
    .A2(_10617_),
    .A3(_10623_),
    .ZN(_10624_));
 BUF_X8 _16457_ (.A(_10577_),
    .Z(_10625_));
 BUF_X8 _16458_ (.A(_10625_),
    .Z(_10626_));
 BUF_X8 _16459_ (.A(_10626_),
    .Z(_10627_));
 BUF_X4 _16460_ (.A(_10627_),
    .Z(_10628_));
 BUF_X4 _16461_ (.A(_10628_),
    .Z(_10629_));
 OR2_X1 _16462_ (.A1(_00141_),
    .A2(_10629_),
    .ZN(_10630_));
 INV_X1 _16463_ (.A(_10583_),
    .ZN(_10631_));
 BUF_X4 _16464_ (.A(_10631_),
    .Z(_10632_));
 OAI21_X1 _16465_ (.A(_10576_),
    .B1(_10630_),
    .B2(_10632_),
    .ZN(_10633_));
 OAI21_X1 _16466_ (.A(_10610_),
    .B1(_10624_),
    .B2(_10633_),
    .ZN(_10634_));
 MUX2_X1 _16467_ (.A(_00159_),
    .B(_00161_),
    .S(_10588_),
    .Z(_10635_));
 MUX2_X1 _16468_ (.A(_00160_),
    .B(_00162_),
    .S(_10588_),
    .Z(_10636_));
 MUX2_X1 _16469_ (.A(_10635_),
    .B(_10636_),
    .S(_10629_),
    .Z(_10637_));
 MUX2_X1 _16470_ (.A(_00143_),
    .B(_00145_),
    .S(_10588_),
    .Z(_10638_));
 MUX2_X1 _16471_ (.A(_00144_),
    .B(_00146_),
    .S(_10588_),
    .Z(_10639_));
 MUX2_X1 _16472_ (.A(_10638_),
    .B(_10639_),
    .S(_10629_),
    .Z(_10640_));
 MUX2_X1 _16473_ (.A(_10637_),
    .B(_10640_),
    .S(_10576_),
    .Z(_10641_));
 OAI221_X2 _16474_ (.A(_10571_),
    .B1(_10605_),
    .B2(_10634_),
    .C1(_10641_),
    .C2(_10610_),
    .ZN(_10642_));
 NOR2_X4 _16475_ (.A1(_10606_),
    .A2(_10567_),
    .ZN(_10643_));
 MUX2_X1 _16476_ (.A(_00163_),
    .B(_00165_),
    .S(_10588_),
    .Z(_10644_));
 MUX2_X1 _16477_ (.A(_00164_),
    .B(_00166_),
    .S(_10621_),
    .Z(_10645_));
 MUX2_X1 _16478_ (.A(_10644_),
    .B(_10645_),
    .S(_10629_),
    .Z(_10646_));
 MUX2_X1 _16479_ (.A(_00147_),
    .B(_00149_),
    .S(_10621_),
    .Z(_10647_));
 MUX2_X1 _16480_ (.A(_00148_),
    .B(_00150_),
    .S(_10621_),
    .Z(_10648_));
 MUX2_X1 _16481_ (.A(_10647_),
    .B(_10648_),
    .S(_10629_),
    .Z(_10649_));
 MUX2_X1 _16482_ (.A(_10646_),
    .B(_10649_),
    .S(_10576_),
    .Z(_10650_));
 NOR2_X2 _16483_ (.A1(_10607_),
    .A2(_10567_),
    .ZN(_10651_));
 MUX2_X1 _16484_ (.A(_00167_),
    .B(_00169_),
    .S(_10601_),
    .Z(_10652_));
 MUX2_X1 _16485_ (.A(_00168_),
    .B(_00170_),
    .S(_10601_),
    .Z(_10653_));
 MUX2_X1 _16486_ (.A(_10652_),
    .B(_10653_),
    .S(_10596_),
    .Z(_10654_));
 MUX2_X1 _16487_ (.A(_00151_),
    .B(_00153_),
    .S(_10601_),
    .Z(_10655_));
 MUX2_X1 _16488_ (.A(_00152_),
    .B(_00154_),
    .S(_10601_),
    .Z(_10656_));
 MUX2_X1 _16489_ (.A(_10655_),
    .B(_10656_),
    .S(_10629_),
    .Z(_10657_));
 MUX2_X1 _16490_ (.A(_10654_),
    .B(_10657_),
    .S(_10576_),
    .Z(_10658_));
 AOI22_X4 _16491_ (.A1(_10643_),
    .A2(_10650_),
    .B1(_10651_),
    .B2(_10658_),
    .ZN(_10659_));
 NAND3_X2 _16492_ (.A1(_10565_),
    .A2(_10642_),
    .A3(_10659_),
    .ZN(_10660_));
 NOR3_X4 _16493_ (.A1(_10292_),
    .A2(_10296_),
    .A3(_10556_),
    .ZN(_10661_));
 AOI22_X4 _16494_ (.A1(_10536_),
    .A2(_10535_),
    .B1(_10661_),
    .B2(_10348_),
    .ZN(_10662_));
 NAND4_X1 _16495_ (.A1(_10341_),
    .A2(_10287_),
    .A3(_10302_),
    .A4(_10330_),
    .ZN(_10663_));
 OAI21_X2 _16496_ (.A(_10663_),
    .B1(_10331_),
    .B2(_10287_),
    .ZN(_10664_));
 AND2_X1 _16497_ (.A1(_10299_),
    .A2(_10513_),
    .ZN(_10665_));
 NAND2_X1 _16498_ (.A1(_10327_),
    .A2(_10312_),
    .ZN(_10666_));
 OAI221_X2 _16499_ (.A(_10555_),
    .B1(_10665_),
    .B2(_10480_),
    .C1(_10384_),
    .C2(_10666_),
    .ZN(_10667_));
 OAI211_X4 _16500_ (.A(_10326_),
    .B(_10662_),
    .C1(_10664_),
    .C2(_10667_),
    .ZN(_10668_));
 AOI21_X4 _16501_ (.A(_10347_),
    .B1(_10555_),
    .B2(_10557_),
    .ZN(_10669_));
 NOR2_X4 _16502_ (.A1(_10344_),
    .A2(_10381_),
    .ZN(_10670_));
 OAI33_X1 _16503_ (.A1(_10666_),
    .A2(_10333_),
    .A3(_10384_),
    .B1(_10340_),
    .B2(_10378_),
    .B3(_10670_),
    .ZN(_10671_));
 OR3_X4 _16504_ (.A1(_10562_),
    .A2(_10669_),
    .A3(_10671_),
    .ZN(_10672_));
 BUF_X8 _16505_ (.A(_10326_),
    .Z(_10673_));
 AOI22_X4 _16506_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(_10668_),
    .B1(_10672_),
    .B2(_10673_),
    .ZN(_10674_));
 CLKBUF_X2 _16507_ (.A(\cs_registers_i.pc_id_i[1] ),
    .Z(_10675_));
 INV_X1 _16508_ (.A(_10675_),
    .ZN(_10676_));
 NAND2_X4 _16509_ (.A1(_10380_),
    .A2(_10346_),
    .ZN(_10677_));
 NOR2_X4 _16510_ (.A1(_10348_),
    .A2(_10677_),
    .ZN(_10678_));
 OR3_X1 _16511_ (.A1(_00183_),
    .A2(_10557_),
    .A3(_10678_),
    .ZN(_10679_));
 MUX2_X1 _16512_ (.A(_10676_),
    .B(_10679_),
    .S(_10668_),
    .Z(_10680_));
 NOR3_X4 _16513_ (.A1(_10562_),
    .A2(_10669_),
    .A3(_10671_),
    .ZN(_10681_));
 NOR2_X4 _16514_ (.A1(_10361_),
    .A2(_10681_),
    .ZN(_10682_));
 BUF_X8 _16515_ (.A(_10682_),
    .Z(_10683_));
 AOI22_X4 _16516_ (.A1(_10660_),
    .A2(_10674_),
    .B1(_10680_),
    .B2(_10683_),
    .ZN(_15845_));
 INV_X1 _16517_ (.A(_15845_),
    .ZN(_15849_));
 BUF_X4 _16518_ (.A(_10430_),
    .Z(_10684_));
 BUF_X4 _16519_ (.A(_10684_),
    .Z(_10685_));
 MUX2_X1 _16520_ (.A(_00208_),
    .B(_00212_),
    .S(_10685_),
    .Z(_10686_));
 MUX2_X1 _16521_ (.A(_00210_),
    .B(_00214_),
    .S(_10685_),
    .Z(_10687_));
 MUX2_X1 _16522_ (.A(_10686_),
    .B(_10687_),
    .S(_10454_),
    .Z(_10688_));
 MUX2_X1 _16523_ (.A(_00192_),
    .B(_00196_),
    .S(_10685_),
    .Z(_10689_));
 MUX2_X1 _16524_ (.A(_00194_),
    .B(_00198_),
    .S(_10685_),
    .Z(_10690_));
 MUX2_X1 _16525_ (.A(_10689_),
    .B(_10690_),
    .S(net357),
    .Z(_10691_));
 MUX2_X1 _16526_ (.A(_10688_),
    .B(_10691_),
    .S(_10473_),
    .Z(_10692_));
 NOR2_X1 _16527_ (.A1(_10466_),
    .A2(_10692_),
    .ZN(_10693_));
 INV_X2 _16528_ (.A(_10412_),
    .ZN(_10694_));
 BUF_X4 _16529_ (.A(_10694_),
    .Z(_10695_));
 BUF_X4 _16530_ (.A(_10695_),
    .Z(_10696_));
 BUF_X4 _16531_ (.A(_10696_),
    .Z(_10697_));
 MUX2_X1 _16532_ (.A(_00209_),
    .B(_00213_),
    .S(_10431_),
    .Z(_10698_));
 MUX2_X1 _16533_ (.A(_00211_),
    .B(_00215_),
    .S(_10685_),
    .Z(_10699_));
 MUX2_X1 _16534_ (.A(_10698_),
    .B(_10699_),
    .S(_10454_),
    .Z(_10700_));
 MUX2_X1 _16535_ (.A(_00193_),
    .B(_00197_),
    .S(_10685_),
    .Z(_10701_));
 MUX2_X1 _16536_ (.A(_00195_),
    .B(_00199_),
    .S(_10685_),
    .Z(_10702_));
 MUX2_X1 _16537_ (.A(_10701_),
    .B(_10702_),
    .S(_10454_),
    .Z(_10703_));
 MUX2_X1 _16538_ (.A(_10700_),
    .B(_10703_),
    .S(_10473_),
    .Z(_10704_));
 NOR2_X1 _16539_ (.A1(_10697_),
    .A2(_10704_),
    .ZN(_10705_));
 NOR3_X2 _16540_ (.A1(_10421_),
    .A2(_10693_),
    .A3(_10705_),
    .ZN(_10706_));
 BUF_X4 _16541_ (.A(_10471_),
    .Z(_10707_));
 BUF_X8 _16542_ (.A(_10707_),
    .Z(_10708_));
 BUF_X4 _16543_ (.A(_10708_),
    .Z(_10709_));
 BUF_X4 _16544_ (.A(_10452_),
    .Z(_10710_));
 MUX2_X1 _16545_ (.A(_00200_),
    .B(_00202_),
    .S(_10710_),
    .Z(_10711_));
 MUX2_X1 _16546_ (.A(_00201_),
    .B(_00203_),
    .S(_10710_),
    .Z(_10712_));
 MUX2_X1 _16547_ (.A(_10711_),
    .B(_10712_),
    .S(_10465_),
    .Z(_10713_));
 NAND2_X1 _16548_ (.A1(_10709_),
    .A2(_10713_),
    .ZN(_10714_));
 NAND2_X4 _16549_ (.A1(_10695_),
    .A2(_10406_),
    .ZN(_10715_));
 BUF_X4 _16550_ (.A(_10715_),
    .Z(_10716_));
 NAND2_X1 _16551_ (.A1(net357),
    .A2(_00187_),
    .ZN(_10717_));
 OAI21_X1 _16552_ (.A(_10717_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B2(net357),
    .ZN(_10718_));
 OAI221_X1 _16553_ (.A(_10474_),
    .B1(_00186_),
    .B2(_10716_),
    .C1(_10718_),
    .C2(_10697_),
    .ZN(_10719_));
 AND3_X1 _16554_ (.A1(_10436_),
    .A2(_10714_),
    .A3(_10719_),
    .ZN(_10720_));
 MUX2_X1 _16555_ (.A(_00204_),
    .B(_00206_),
    .S(_10406_),
    .Z(_10721_));
 MUX2_X1 _16556_ (.A(_00205_),
    .B(_00207_),
    .S(_10406_),
    .Z(_10722_));
 MUX2_X1 _16557_ (.A(_10721_),
    .B(_10722_),
    .S(_10414_),
    .Z(_10723_));
 MUX2_X1 _16558_ (.A(_00188_),
    .B(_00190_),
    .S(_10406_),
    .Z(_10724_));
 MUX2_X1 _16559_ (.A(_00189_),
    .B(_00191_),
    .S(_10406_),
    .Z(_10725_));
 MUX2_X1 _16560_ (.A(_10724_),
    .B(_10725_),
    .S(_10414_),
    .Z(_10726_));
 MUX2_X1 _16561_ (.A(_10723_),
    .B(_10726_),
    .S(_10473_),
    .Z(_10727_));
 NOR2_X1 _16562_ (.A1(_10436_),
    .A2(_10727_),
    .ZN(_10728_));
 NOR3_X2 _16563_ (.A1(_10468_),
    .A2(_10720_),
    .A3(_10728_),
    .ZN(_10729_));
 NOR3_X4 _16564_ (.A1(_10317_),
    .A2(_10706_),
    .A3(_10729_),
    .ZN(_10730_));
 INV_X1 _16565_ (.A(_00216_),
    .ZN(_10731_));
 AOI211_X2 _16566_ (.A(_10731_),
    .B(_10360_),
    .C1(_10371_),
    .C2(_10375_),
    .ZN(_10732_));
 NAND3_X1 _16567_ (.A1(_10317_),
    .A2(_10389_),
    .A3(_10386_),
    .ZN(_10733_));
 OAI21_X1 _16568_ (.A(_10673_),
    .B1(_10374_),
    .B2(net18),
    .ZN(_10734_));
 AOI211_X2 _16569_ (.A(_10732_),
    .B(_10733_),
    .C1(_10734_),
    .C2(_10697_),
    .ZN(_10735_));
 OAI21_X4 _16570_ (.A(_10673_),
    .B1(_10735_),
    .B2(_10730_),
    .ZN(_10736_));
 INV_X1 _16571_ (.A(_10736_),
    .ZN(_10737_));
 BUF_X4 _16572_ (.A(_10737_),
    .Z(_10738_));
 BUF_X4 _16573_ (.A(_10738_),
    .Z(_15841_));
 BUF_X8 _16574_ (.A(_10736_),
    .Z(_10739_));
 BUF_X1 rebuffer7 (.A(_11500_),
    .Z(net278));
 BUF_X4 _16576_ (.A(_10739_),
    .Z(_15835_));
 BUF_X8 _16577_ (.A(_10361_),
    .Z(_10741_));
 NAND2_X2 _16578_ (.A1(_10522_),
    .A2(_10670_),
    .ZN(_10742_));
 NAND2_X1 _16579_ (.A1(_10661_),
    .A2(_10742_),
    .ZN(_10743_));
 BUF_X4 _16580_ (.A(_10743_),
    .Z(_10744_));
 NOR4_X1 _16581_ (.A1(_00184_),
    .A2(_10741_),
    .A3(_10681_),
    .A4(_10744_),
    .ZN(_10745_));
 NAND2_X2 _16582_ (.A1(_10326_),
    .A2(_10672_),
    .ZN(_10746_));
 BUF_X4 _16583_ (.A(_10746_),
    .Z(_10747_));
 AOI21_X2 _16584_ (.A(_10745_),
    .B1(_10747_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .ZN(_10748_));
 BUF_X8 _16585_ (.A(_10572_),
    .Z(_10749_));
 BUF_X8 _16586_ (.A(_10749_),
    .Z(_10750_));
 BUF_X4 _16587_ (.A(_10606_),
    .Z(_10751_));
 BUF_X8 _16588_ (.A(_10751_),
    .Z(_10752_));
 MUX2_X1 _16589_ (.A(_00188_),
    .B(_00190_),
    .S(_10589_),
    .Z(_10753_));
 MUX2_X1 _16590_ (.A(_00189_),
    .B(_00191_),
    .S(_10589_),
    .Z(_10754_));
 MUX2_X1 _16591_ (.A(_10753_),
    .B(_10754_),
    .S(_10597_),
    .Z(_10755_));
 NAND2_X1 _16592_ (.A1(_10752_),
    .A2(_10755_),
    .ZN(_10756_));
 NAND2_X4 _16593_ (.A1(_10580_),
    .A2(_10601_),
    .ZN(_10757_));
 BUF_X4 _16594_ (.A(_10757_),
    .Z(_10758_));
 BUF_X8 _16595_ (.A(_10622_),
    .Z(_10759_));
 NAND2_X1 _16596_ (.A1(_10759_),
    .A2(_00187_),
    .ZN(_10760_));
 OAI21_X1 _16597_ (.A(_10760_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B2(_10759_),
    .ZN(_10761_));
 OAI221_X1 _16598_ (.A(_10610_),
    .B1(_00186_),
    .B2(_10758_),
    .C1(_10761_),
    .C2(_10582_),
    .ZN(_10762_));
 NAND3_X1 _16599_ (.A1(_10571_),
    .A2(_10756_),
    .A3(_10762_),
    .ZN(_10763_));
 BUF_X8 _16600_ (.A(_10566_),
    .Z(_10764_));
 BUF_X4 _16601_ (.A(_10764_),
    .Z(_10765_));
 BUF_X4 _16602_ (.A(_10765_),
    .Z(_10766_));
 BUF_X4 _16603_ (.A(_10766_),
    .Z(_10767_));
 MUX2_X1 _16604_ (.A(_00194_),
    .B(_00198_),
    .S(_10751_),
    .Z(_10768_));
 MUX2_X1 _16605_ (.A(_00195_),
    .B(_00199_),
    .S(_10751_),
    .Z(_10769_));
 MUX2_X1 _16606_ (.A(_10768_),
    .B(_10769_),
    .S(_10597_),
    .Z(_10770_));
 NAND2_X1 _16607_ (.A1(_10759_),
    .A2(_10770_),
    .ZN(_10771_));
 MUX2_X1 _16608_ (.A(_00192_),
    .B(_00196_),
    .S(_10751_),
    .Z(_10772_));
 MUX2_X1 _16609_ (.A(_00193_),
    .B(_00197_),
    .S(_10751_),
    .Z(_10773_));
 MUX2_X1 _16610_ (.A(_10772_),
    .B(_10773_),
    .S(_10597_),
    .Z(_10774_));
 NAND2_X1 _16611_ (.A1(_10632_),
    .A2(_10774_),
    .ZN(_10775_));
 NAND3_X1 _16612_ (.A1(_10767_),
    .A2(_10771_),
    .A3(_10775_),
    .ZN(_10776_));
 AOI21_X2 _16613_ (.A(_10750_),
    .B1(_10763_),
    .B2(_10776_),
    .ZN(_10777_));
 NOR2_X4 _16614_ (.A1(_10607_),
    .A2(_10764_),
    .ZN(_10778_));
 MUX2_X1 _16615_ (.A(_00204_),
    .B(_00206_),
    .S(_10589_),
    .Z(_10779_));
 MUX2_X1 _16616_ (.A(_00205_),
    .B(_00207_),
    .S(_10589_),
    .Z(_10780_));
 MUX2_X1 _16617_ (.A(_10779_),
    .B(_10780_),
    .S(_10597_),
    .Z(_10781_));
 NAND2_X1 _16618_ (.A1(_10778_),
    .A2(_10781_),
    .ZN(_10782_));
 BUF_X8 _16619_ (.A(_10574_),
    .Z(_10783_));
 NOR3_X4 _16620_ (.A1(_10585_),
    .A2(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .A3(_10764_),
    .ZN(_10784_));
 BUF_X8 _16621_ (.A(_10784_),
    .Z(_10785_));
 BUF_X4 _16622_ (.A(_10625_),
    .Z(_10786_));
 BUF_X4 _16623_ (.A(_10786_),
    .Z(_10787_));
 BUF_X4 _16624_ (.A(_10787_),
    .Z(_10788_));
 MUX2_X1 _16625_ (.A(_00200_),
    .B(_00201_),
    .S(_10788_),
    .Z(_10789_));
 BUF_X4 _16626_ (.A(_10583_),
    .Z(_10790_));
 BUF_X4 _16627_ (.A(_10790_),
    .Z(_10791_));
 NOR2_X2 _16628_ (.A1(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .A2(_10566_),
    .ZN(_10792_));
 AND2_X1 _16629_ (.A1(_10791_),
    .A2(_10792_),
    .ZN(_10793_));
 BUF_X8 _16630_ (.A(_10793_),
    .Z(_10794_));
 BUF_X8 _16631_ (.A(_10625_),
    .Z(_10795_));
 BUF_X4 _16632_ (.A(_10795_),
    .Z(_10796_));
 BUF_X8 _16633_ (.A(_10796_),
    .Z(_10797_));
 MUX2_X1 _16634_ (.A(_00202_),
    .B(_00203_),
    .S(_10797_),
    .Z(_10798_));
 AOI221_X2 _16635_ (.A(_10783_),
    .B1(_10785_),
    .B2(_10789_),
    .C1(_10794_),
    .C2(_10798_),
    .ZN(_10799_));
 MUX2_X1 _16636_ (.A(_00214_),
    .B(_00215_),
    .S(_10797_),
    .Z(_10800_));
 AOI21_X1 _16637_ (.A(_10609_),
    .B1(_10800_),
    .B2(_10616_),
    .ZN(_10801_));
 MUX2_X1 _16638_ (.A(_00210_),
    .B(_00211_),
    .S(_10788_),
    .Z(_10802_));
 AOI21_X1 _16639_ (.A(_10752_),
    .B1(_10802_),
    .B2(_10616_),
    .ZN(_10803_));
 OAI21_X1 _16640_ (.A(_10759_),
    .B1(_10801_),
    .B2(_10803_),
    .ZN(_10804_));
 NAND2_X1 _16641_ (.A1(_10582_),
    .A2(_00208_),
    .ZN(_10805_));
 NAND2_X1 _16642_ (.A1(_10597_),
    .A2(_00209_),
    .ZN(_10806_));
 NAND3_X1 _16643_ (.A1(_10803_),
    .A2(_10805_),
    .A3(_10806_),
    .ZN(_10807_));
 NAND2_X1 _16644_ (.A1(_10582_),
    .A2(_00212_),
    .ZN(_10808_));
 NAND2_X1 _16645_ (.A1(_10597_),
    .A2(_00213_),
    .ZN(_10809_));
 NAND3_X1 _16646_ (.A1(_10801_),
    .A2(_10808_),
    .A3(_10809_),
    .ZN(_10810_));
 NAND4_X1 _16647_ (.A1(_10767_),
    .A2(_10804_),
    .A3(_10807_),
    .A4(_10810_),
    .ZN(_10811_));
 AND3_X1 _16648_ (.A1(_10782_),
    .A2(_10799_),
    .A3(_10811_),
    .ZN(_10812_));
 NOR2_X4 _16649_ (.A1(_10812_),
    .A2(_10777_),
    .ZN(_10813_));
 NAND2_X4 _16650_ (.A1(_10563_),
    .A2(_10746_),
    .ZN(_10814_));
 OAI22_X4 _16651_ (.A1(_10565_),
    .A2(_10748_),
    .B1(_10813_),
    .B2(_10814_),
    .ZN(_15842_));
 INV_X2 _16652_ (.A(_15842_),
    .ZN(_15838_));
 BUF_X4 _16653_ (.A(_15372_),
    .Z(_10815_));
 XOR2_X2 _16654_ (.A(_14067_),
    .B(_10815_),
    .Z(\alu_adder_result_ex[1] ));
 INV_X4 _16655_ (.A(net15),
    .ZN(_16090_));
 AOI21_X4 _16656_ (.A(_10668_),
    .B1(_10672_),
    .B2(_10673_),
    .ZN(_10816_));
 MUX2_X1 _16657_ (.A(_00224_),
    .B(_00226_),
    .S(_10619_),
    .Z(_10817_));
 MUX2_X1 _16658_ (.A(_00225_),
    .B(_00227_),
    .S(_10619_),
    .Z(_10818_));
 MUX2_X1 _16659_ (.A(_10817_),
    .B(_10818_),
    .S(_10796_),
    .Z(_10819_));
 INV_X1 _16660_ (.A(_00218_),
    .ZN(_10820_));
 NOR2_X4 _16661_ (.A1(_10577_),
    .A2(_10631_),
    .ZN(_10821_));
 BUF_X4 _16662_ (.A(_10821_),
    .Z(_10822_));
 BUF_X4 _16663_ (.A(_10599_),
    .Z(_10823_));
 NOR2_X1 _16664_ (.A1(_10823_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .ZN(_10824_));
 AOI21_X1 _16665_ (.A(_10824_),
    .B1(_00219_),
    .B2(_10614_),
    .ZN(_10825_));
 AOI22_X1 _16666_ (.A1(_10820_),
    .A2(_10822_),
    .B1(_10825_),
    .B2(_10595_),
    .ZN(_10826_));
 BUF_X4 _16667_ (.A(_10567_),
    .Z(_10827_));
 BUF_X4 _16668_ (.A(_10827_),
    .Z(_10828_));
 MUX2_X1 _16669_ (.A(_10819_),
    .B(_10826_),
    .S(_10828_),
    .Z(_10829_));
 NAND2_X1 _16670_ (.A1(_10607_),
    .A2(_10573_),
    .ZN(_10830_));
 BUF_X4 _16671_ (.A(_10830_),
    .Z(_10831_));
 BUF_X4 _16672_ (.A(_10606_),
    .Z(_10832_));
 BUF_X4 _16673_ (.A(_10592_),
    .Z(_10833_));
 MUX2_X1 _16674_ (.A(_00242_),
    .B(_00243_),
    .S(_10833_),
    .Z(_10834_));
 MUX2_X1 _16675_ (.A(_00240_),
    .B(_00241_),
    .S(_10833_),
    .Z(_10835_));
 MUX2_X1 _16676_ (.A(_10834_),
    .B(_10835_),
    .S(_10632_),
    .Z(_10836_));
 NOR2_X1 _16677_ (.A1(_10832_),
    .A2(_10836_),
    .ZN(_10837_));
 NAND2_X1 _16678_ (.A1(_10601_),
    .A2(_10606_),
    .ZN(_10838_));
 BUF_X4 _16679_ (.A(_10592_),
    .Z(_10839_));
 BUF_X1 rebuffer88 (.A(net358),
    .Z(net359));
 MUX2_X1 _16681_ (.A(_00246_),
    .B(_00247_),
    .S(_10839_),
    .Z(_10841_));
 NAND2_X1 _16682_ (.A1(_10632_),
    .A2(_10606_),
    .ZN(_10842_));
 BUF_X4 _16683_ (.A(_10625_),
    .Z(_10843_));
 MUX2_X1 _16684_ (.A(_00244_),
    .B(_00245_),
    .S(_10843_),
    .Z(_10844_));
 OAI22_X1 _16685_ (.A1(_10838_),
    .A2(_10841_),
    .B1(_10842_),
    .B2(_10844_),
    .ZN(_10845_));
 NOR3_X1 _16686_ (.A1(_10570_),
    .A2(_10837_),
    .A3(_10845_),
    .ZN(_10846_));
 MUX2_X1 _16687_ (.A(_00236_),
    .B(_00238_),
    .S(_10619_),
    .Z(_10847_));
 MUX2_X1 _16688_ (.A(_00237_),
    .B(_00239_),
    .S(_10619_),
    .Z(_10848_));
 MUX2_X1 _16689_ (.A(_10847_),
    .B(_10848_),
    .S(_10787_),
    .Z(_10849_));
 NAND2_X1 _16690_ (.A1(_10778_),
    .A2(_10849_),
    .ZN(_10850_));
 MUX2_X1 _16691_ (.A(_00232_),
    .B(_00233_),
    .S(_10625_),
    .Z(_10851_));
 MUX2_X1 _16692_ (.A(_00234_),
    .B(_00235_),
    .S(_10593_),
    .Z(_10852_));
 AOI221_X1 _16693_ (.A(_10573_),
    .B1(_10784_),
    .B2(_10851_),
    .C1(_10852_),
    .C2(_10794_),
    .ZN(_10853_));
 NAND2_X1 _16694_ (.A1(_10850_),
    .A2(_10853_),
    .ZN(_10854_));
 NAND2_X4 _16695_ (.A1(_10606_),
    .A2(_10573_),
    .ZN(_10855_));
 BUF_X8 _16696_ (.A(_10583_),
    .Z(_10856_));
 BUF_X8 _16697_ (.A(_10856_),
    .Z(_10857_));
 BUF_X4 _16698_ (.A(_10857_),
    .Z(_10858_));
 MUX2_X1 _16699_ (.A(_00228_),
    .B(_00230_),
    .S(_10858_),
    .Z(_10859_));
 MUX2_X1 _16700_ (.A(_00229_),
    .B(_00231_),
    .S(_10858_),
    .Z(_10860_));
 BUF_X8 _16701_ (.A(_10592_),
    .Z(_10861_));
 BUF_X8 _16702_ (.A(_10861_),
    .Z(_10862_));
 MUX2_X1 _16703_ (.A(_10859_),
    .B(_10860_),
    .S(_10862_),
    .Z(_10863_));
 MUX2_X1 _16704_ (.A(_00220_),
    .B(_00222_),
    .S(_10858_),
    .Z(_10864_));
 MUX2_X1 _16705_ (.A(_00221_),
    .B(_00223_),
    .S(_10858_),
    .Z(_10865_));
 MUX2_X1 _16706_ (.A(_10864_),
    .B(_10865_),
    .S(_10594_),
    .Z(_10866_));
 MUX2_X1 _16707_ (.A(_10863_),
    .B(_10866_),
    .S(_10569_),
    .Z(_10867_));
 OAI222_X2 _16708_ (.A1(_10829_),
    .A2(_10831_),
    .B1(_10846_),
    .B2(_10854_),
    .C1(_10855_),
    .C2(_10867_),
    .ZN(_10868_));
 AND2_X1 _16709_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_10563_),
    .ZN(_10869_));
 BUF_X4 _16710_ (.A(_10682_),
    .Z(_10870_));
 AOI222_X2 _16711_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(_10741_),
    .B1(_10816_),
    .B2(_10868_),
    .C1(_10869_),
    .C2(_10870_),
    .ZN(_15936_));
 NAND2_X1 _16712_ (.A1(_10661_),
    .A2(_10670_),
    .ZN(_10871_));
 BUF_X4 _16713_ (.A(_10707_),
    .Z(_10872_));
 BUF_X4 _16714_ (.A(_10507_),
    .Z(_10873_));
 BUF_X4 _16715_ (.A(\id_stage_i.controller_i.instr_i[26] ),
    .Z(_10874_));
 NOR4_X2 _16716_ (.A1(_10872_),
    .A2(_10873_),
    .A3(_10500_),
    .A4(_10874_),
    .ZN(_10875_));
 NAND2_X4 _16717_ (.A1(_10540_),
    .A2(_10875_),
    .ZN(_10876_));
 INV_X1 _16718_ (.A(_10502_),
    .ZN(_10877_));
 NAND2_X1 _16719_ (.A1(net305),
    .A2(_10877_),
    .ZN(_10878_));
 BUF_X4 _16720_ (.A(_10412_),
    .Z(_10879_));
 NAND2_X4 _16721_ (.A1(_10879_),
    .A2(_10337_),
    .ZN(_10880_));
 NAND2_X4 _16722_ (.A1(_10685_),
    .A2(_10421_),
    .ZN(_10881_));
 NOR4_X4 _16723_ (.A1(_10876_),
    .A2(_10878_),
    .A3(_10880_),
    .A4(_10881_),
    .ZN(_10882_));
 OR2_X2 _16724_ (.A1(_10509_),
    .A2(_10498_),
    .ZN(_10883_));
 OR3_X1 _16725_ (.A1(_10500_),
    .A2(_10874_),
    .A3(_10883_),
    .ZN(_10884_));
 NAND2_X2 _16726_ (.A1(net305),
    .A2(_10502_),
    .ZN(_10885_));
 OR3_X4 _16727_ (.A1(_10413_),
    .A2(_10337_),
    .A3(_10885_),
    .ZN(_10886_));
 NAND2_X2 _16728_ (.A1(_10510_),
    .A2(_10498_),
    .ZN(_10887_));
 INV_X2 _16729_ (.A(_10874_),
    .ZN(_10888_));
 NAND4_X4 _16730_ (.A1(_10708_),
    .A2(_10873_),
    .A3(_10500_),
    .A4(_10888_),
    .ZN(_10889_));
 OAI33_X1 _16731_ (.A1(_10709_),
    .A2(_10873_),
    .A3(_10884_),
    .B1(_10886_),
    .B2(_10887_),
    .B3(_10889_),
    .ZN(_10890_));
 NAND2_X4 _16732_ (.A1(_10435_),
    .A2(_10420_),
    .ZN(_10891_));
 OR3_X2 _16733_ (.A1(net397),
    .A2(net305),
    .A3(_10502_),
    .ZN(_10892_));
 AOI21_X1 _16734_ (.A(_10891_),
    .B1(_10886_),
    .B2(_10892_),
    .ZN(_10893_));
 AOI211_X2 _16735_ (.A(_10871_),
    .B(_10882_),
    .C1(_10890_),
    .C2(_10893_),
    .ZN(_10894_));
 NOR4_X4 _16736_ (.A1(_10289_),
    .A2(_10292_),
    .A3(_10296_),
    .A4(_10307_),
    .ZN(_10895_));
 NOR2_X1 _16737_ (.A1(_10310_),
    .A2(_00175_),
    .ZN(_10896_));
 AOI21_X2 _16738_ (.A(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .B1(_10895_),
    .B2(_10896_),
    .ZN(_10897_));
 NAND3_X4 _16739_ (.A1(_10580_),
    .A2(_00180_),
    .A3(_10784_),
    .ZN(_10898_));
 CLKBUF_X3 _16740_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Z(_10899_));
 INV_X1 _16741_ (.A(_10899_),
    .ZN(_10900_));
 INV_X2 _16742_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .ZN(_10901_));
 BUF_X4 _16743_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .Z(_10902_));
 BUF_X4 _16744_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .Z(_10903_));
 NOR3_X4 _16745_ (.A1(_10394_),
    .A2(_10902_),
    .A3(_10903_),
    .ZN(_10904_));
 NAND4_X1 _16746_ (.A1(_10522_),
    .A2(_10900_),
    .A3(_10901_),
    .A4(_10904_),
    .ZN(_10905_));
 NOR2_X1 _16747_ (.A1(_10898_),
    .A2(_10905_),
    .ZN(_10906_));
 OAI21_X1 _16748_ (.A(_10346_),
    .B1(_10402_),
    .B2(_10287_),
    .ZN(_10907_));
 AOI22_X1 _16749_ (.A1(_10287_),
    .A2(_10348_),
    .B1(_10907_),
    .B2(_10344_),
    .ZN(_10908_));
 BUF_X4 _16750_ (.A(_10315_),
    .Z(_10909_));
 OAI221_X2 _16751_ (.A(_10897_),
    .B1(_10871_),
    .B2(_10906_),
    .C1(_10908_),
    .C2(_10909_),
    .ZN(_10910_));
 OR4_X4 _16752_ (.A1(_10296_),
    .A2(_10292_),
    .A3(_10298_),
    .A4(_10513_),
    .ZN(_10911_));
 BUF_X16 _16753_ (.A(_10911_),
    .Z(_10912_));
 AND2_X1 _16754_ (.A1(_10511_),
    .A2(_10543_),
    .ZN(_10913_));
 XNOR2_X1 _16755_ (.A(_10310_),
    .B(_10381_),
    .ZN(_10914_));
 NAND2_X1 _16756_ (.A1(_10508_),
    .A2(_10914_),
    .ZN(_10915_));
 OR4_X2 _16757_ (.A1(_10500_),
    .A2(_10874_),
    .A3(_10501_),
    .A4(_10502_),
    .ZN(_10916_));
 NOR2_X4 _16758_ (.A1(_10916_),
    .A2(_10883_),
    .ZN(_10917_));
 AOI221_X2 _16759_ (.A(_10912_),
    .B1(_10913_),
    .B2(_10914_),
    .C1(_10915_),
    .C2(_10917_),
    .ZN(_10918_));
 OR4_X4 _16760_ (.A1(_10744_),
    .A2(_10894_),
    .A3(_10910_),
    .A4(_10918_),
    .ZN(_10919_));
 BUF_X4 _16761_ (.A(_10919_),
    .Z(_10920_));
 NOR2_X2 _16762_ (.A1(_15835_),
    .A2(_10920_),
    .ZN(_15511_));
 INV_X1 _16763_ (.A(_15511_),
    .ZN(_15514_));
 NOR4_X4 _16764_ (.A1(_10744_),
    .A2(_10894_),
    .A3(_10910_),
    .A4(_10918_),
    .ZN(_10921_));
 BUF_X4 _16765_ (.A(_10921_),
    .Z(_10922_));
 NAND2_X2 _16766_ (.A1(_15846_),
    .A2(_10922_),
    .ZN(_15510_));
 INV_X1 _16767_ (.A(_15510_),
    .ZN(_15517_));
 NAND2_X2 _16768_ (.A1(_10326_),
    .A2(_10316_),
    .ZN(_10923_));
 NAND3_X1 _16769_ (.A1(_10432_),
    .A2(_10371_),
    .A3(_10375_),
    .ZN(_10924_));
 OAI21_X1 _16770_ (.A(_00278_),
    .B1(_10361_),
    .B2(_10354_),
    .ZN(_10925_));
 NOR2_X4 _16771_ (.A1(_10374_),
    .A2(net19),
    .ZN(_10926_));
 OAI21_X1 _16772_ (.A(_10924_),
    .B1(_10925_),
    .B2(_10926_),
    .ZN(_10927_));
 NAND2_X4 _16773_ (.A1(_10330_),
    .A2(_10385_),
    .ZN(_10928_));
 NAND2_X1 _16774_ (.A1(_10326_),
    .A2(_10928_),
    .ZN(_10929_));
 OAI21_X2 _16775_ (.A(_10389_),
    .B1(_10374_),
    .B2(net20),
    .ZN(_10930_));
 NAND3_X2 _16776_ (.A1(_10334_),
    .A2(_10371_),
    .A3(_10375_),
    .ZN(_10931_));
 AOI21_X2 _16777_ (.A(_10929_),
    .B1(_10930_),
    .B2(_10931_),
    .ZN(_10932_));
 AOI221_X2 _16778_ (.A(_10923_),
    .B1(_10927_),
    .B2(_10389_),
    .C1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C2(_10932_),
    .ZN(_10933_));
 BUF_X8 _16779_ (.A(_10933_),
    .Z(_10934_));
 NOR2_X1 _16780_ (.A1(_10435_),
    .A2(_10451_),
    .ZN(_10935_));
 MUX2_X1 _16781_ (.A(_00266_),
    .B(_00268_),
    .S(_10409_),
    .Z(_10936_));
 MUX2_X1 _16782_ (.A(_00267_),
    .B(_00269_),
    .S(_10409_),
    .Z(_10937_));
 MUX2_X1 _16783_ (.A(_10936_),
    .B(_10937_),
    .S(_10413_),
    .Z(_10938_));
 MUX2_X1 _16784_ (.A(_00250_),
    .B(_00252_),
    .S(_10409_),
    .Z(_10939_));
 MUX2_X1 _16785_ (.A(_00251_),
    .B(_00253_),
    .S(_10409_),
    .Z(_10940_));
 BUF_X4 _16786_ (.A(_10879_),
    .Z(_10941_));
 MUX2_X1 _16787_ (.A(_10939_),
    .B(_10940_),
    .S(_10941_),
    .Z(_10942_));
 MUX2_X1 _16788_ (.A(_10938_),
    .B(_10942_),
    .S(_10473_),
    .Z(_10943_));
 AND2_X2 _16789_ (.A1(_10419_),
    .A2(_10471_),
    .ZN(_10944_));
 MUX2_X1 _16790_ (.A(_00271_),
    .B(_00275_),
    .S(_10434_),
    .Z(_10945_));
 MUX2_X1 _16791_ (.A(_00273_),
    .B(_00277_),
    .S(_10434_),
    .Z(_10946_));
 MUX2_X1 _16792_ (.A(_10945_),
    .B(_10946_),
    .S(_10453_),
    .Z(_10947_));
 MUX2_X1 _16793_ (.A(_00270_),
    .B(_00274_),
    .S(_10434_),
    .Z(_10948_));
 MUX2_X1 _16794_ (.A(_00272_),
    .B(_00276_),
    .S(_10434_),
    .Z(_10949_));
 MUX2_X1 _16795_ (.A(_10948_),
    .B(_10949_),
    .S(_10453_),
    .Z(_10950_));
 MUX2_X1 _16796_ (.A(_10947_),
    .B(_10950_),
    .S(_10696_),
    .Z(_10951_));
 AOI22_X2 _16797_ (.A1(_10935_),
    .A2(_10943_),
    .B1(_10944_),
    .B2(_10951_),
    .ZN(_10952_));
 MUX2_X1 _16798_ (.A(_00255_),
    .B(_00257_),
    .S(_10453_),
    .Z(_10953_));
 NOR2_X1 _16799_ (.A1(_10432_),
    .A2(_10953_),
    .ZN(_10954_));
 MUX2_X1 _16800_ (.A(_00259_),
    .B(_00261_),
    .S(_10410_),
    .Z(_10955_));
 NOR2_X1 _16801_ (.A1(_10435_),
    .A2(_10955_),
    .ZN(_10956_));
 OAI21_X1 _16802_ (.A(_10444_),
    .B1(_10954_),
    .B2(_10956_),
    .ZN(_10957_));
 MUX2_X1 _16803_ (.A(_00258_),
    .B(_00260_),
    .S(_10410_),
    .Z(_10958_));
 MUX2_X1 _16804_ (.A(_00254_),
    .B(_00256_),
    .S(_10410_),
    .Z(_10959_));
 MUX2_X1 _16805_ (.A(_10958_),
    .B(_10959_),
    .S(_10435_),
    .Z(_10960_));
 OAI21_X1 _16806_ (.A(_10957_),
    .B1(_10960_),
    .B2(_10466_),
    .ZN(_10961_));
 NAND2_X4 _16807_ (.A1(_10419_),
    .A2(_10472_),
    .ZN(_10962_));
 INV_X1 _16808_ (.A(_00248_),
    .ZN(_10963_));
 NOR2_X4 _16809_ (.A1(_10412_),
    .A2(_10336_),
    .ZN(_10964_));
 NOR2_X1 _16810_ (.A1(_10438_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .ZN(_10965_));
 AOI21_X1 _16811_ (.A(_10965_),
    .B1(_00249_),
    .B2(_10710_),
    .ZN(_10966_));
 AOI221_X2 _16812_ (.A(_10708_),
    .B1(_10963_),
    .B2(_10964_),
    .C1(_10966_),
    .C2(_10443_),
    .ZN(_10967_));
 MUX2_X1 _16813_ (.A(_00262_),
    .B(_00264_),
    .S(_10710_),
    .Z(_10968_));
 MUX2_X1 _16814_ (.A(_00263_),
    .B(_00265_),
    .S(_10710_),
    .Z(_10969_));
 MUX2_X1 _16815_ (.A(_10968_),
    .B(_10969_),
    .S(_10465_),
    .Z(_10970_));
 AOI21_X1 _16816_ (.A(_10967_),
    .B1(_10970_),
    .B2(_10709_),
    .ZN(_10971_));
 OAI221_X2 _16817_ (.A(_10952_),
    .B1(_10961_),
    .B2(_10962_),
    .C1(_10891_),
    .C2(_10971_),
    .ZN(_10972_));
 INV_X4 _16818_ (.A(_10972_),
    .ZN(_10973_));
 NAND2_X4 _16819_ (.A1(_10673_),
    .A2(_10403_),
    .ZN(_10974_));
 NOR2_X4 _16820_ (.A1(_10973_),
    .A2(_10974_),
    .ZN(_10975_));
 NOR2_X4 _16821_ (.A1(_10934_),
    .A2(_10975_),
    .ZN(_15853_));
 INV_X2 _16822_ (.A(_15853_),
    .ZN(_15857_));
 NOR2_X4 _16823_ (.A1(_10360_),
    .A2(_10316_),
    .ZN(_10976_));
 NAND2_X4 _16824_ (.A1(_10442_),
    .A2(_10438_),
    .ZN(_10977_));
 BUF_X4 _16825_ (.A(_10430_),
    .Z(_10978_));
 MUX2_X1 _16826_ (.A(_00304_),
    .B(_00308_),
    .S(_10978_),
    .Z(_10979_));
 OR2_X4 _16827_ (.A1(_10879_),
    .A2(net401),
    .ZN(_10980_));
 MUX2_X1 _16828_ (.A(_00301_),
    .B(_00305_),
    .S(_10684_),
    .Z(_10981_));
 MUX2_X1 _16829_ (.A(_00302_),
    .B(_00306_),
    .S(_10684_),
    .Z(_10982_));
 OAI222_X2 _16830_ (.A1(_10977_),
    .A2(_10979_),
    .B1(_10980_),
    .B2(_10981_),
    .C1(_10982_),
    .C2(_10880_),
    .ZN(_10983_));
 BUF_X4 _16831_ (.A(_10430_),
    .Z(_10984_));
 MUX2_X1 _16832_ (.A(_00303_),
    .B(_00307_),
    .S(_10984_),
    .Z(_10985_));
 OAI21_X1 _16833_ (.A(_10944_),
    .B1(_10985_),
    .B2(_10715_),
    .ZN(_10986_));
 OR2_X1 _16834_ (.A1(_10983_),
    .A2(_10986_),
    .ZN(_10987_));
 NOR2_X4 _16835_ (.A1(_10709_),
    .A2(_10881_),
    .ZN(_10988_));
 MUX2_X1 _16836_ (.A(_00281_),
    .B(_00283_),
    .S(_10405_),
    .Z(_10989_));
 MUX2_X1 _16837_ (.A(_00282_),
    .B(_00284_),
    .S(_10405_),
    .Z(_10990_));
 MUX2_X1 _16838_ (.A(_10989_),
    .B(_10990_),
    .S(_10413_),
    .Z(_10991_));
 MUX2_X1 _16839_ (.A(_00293_),
    .B(_00295_),
    .S(_10405_),
    .Z(_10992_));
 MUX2_X1 _16840_ (.A(_00294_),
    .B(_00296_),
    .S(_10405_),
    .Z(_10993_));
 MUX2_X1 _16841_ (.A(_10992_),
    .B(_10993_),
    .S(_10442_),
    .Z(_10994_));
 NOR2_X4 _16842_ (.A1(_10472_),
    .A2(_10891_),
    .ZN(_10995_));
 AOI22_X1 _16843_ (.A1(_10988_),
    .A2(_10991_),
    .B1(_10994_),
    .B2(_10995_),
    .ZN(_10996_));
 NOR2_X4 _16844_ (.A1(_10430_),
    .A2(_10419_),
    .ZN(_10997_));
 NAND2_X4 _16845_ (.A1(_10472_),
    .A2(_10997_),
    .ZN(_10998_));
 NOR2_X1 _16846_ (.A1(_10408_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .ZN(_10999_));
 AOI21_X1 _16847_ (.A(_10999_),
    .B1(_00280_),
    .B2(_10437_),
    .ZN(_11000_));
 INV_X1 _16848_ (.A(_00279_),
    .ZN(_11001_));
 AOI221_X2 _16849_ (.A(_10998_),
    .B1(_11000_),
    .B2(_10412_),
    .C1(_11001_),
    .C2(_10964_),
    .ZN(_11002_));
 MUX2_X1 _16850_ (.A(_00297_),
    .B(_00299_),
    .S(_10452_),
    .Z(_11003_));
 MUX2_X1 _16851_ (.A(_00298_),
    .B(_00300_),
    .S(_10452_),
    .Z(_11004_));
 MUX2_X1 _16852_ (.A(_11003_),
    .B(_11004_),
    .S(_10941_),
    .Z(_11005_));
 NOR2_X4 _16853_ (.A1(_10472_),
    .A2(_10881_),
    .ZN(_11006_));
 AOI21_X1 _16854_ (.A(_11002_),
    .B1(_11005_),
    .B2(_11006_),
    .ZN(_11007_));
 NOR2_X1 _16855_ (.A1(_10465_),
    .A2(_10962_),
    .ZN(_11008_));
 MUX2_X1 _16856_ (.A(_00285_),
    .B(_00289_),
    .S(_10684_),
    .Z(_11009_));
 MUX2_X1 _16857_ (.A(_00287_),
    .B(_00291_),
    .S(_10684_),
    .Z(_11010_));
 MUX2_X1 _16858_ (.A(_11009_),
    .B(_11010_),
    .S(_10710_),
    .Z(_11011_));
 MUX2_X1 _16859_ (.A(_00286_),
    .B(_00290_),
    .S(_10434_),
    .Z(_11012_));
 MUX2_X1 _16860_ (.A(_00288_),
    .B(_00292_),
    .S(_10434_),
    .Z(_11013_));
 MUX2_X1 _16861_ (.A(_11012_),
    .B(_11013_),
    .S(_10453_),
    .Z(_11014_));
 NAND2_X2 _16862_ (.A1(_10413_),
    .A2(_10451_),
    .ZN(_11015_));
 NOR2_X1 _16863_ (.A1(_10708_),
    .A2(_11015_),
    .ZN(_11016_));
 AOI22_X1 _16864_ (.A1(_11008_),
    .A2(_11011_),
    .B1(_11014_),
    .B2(_11016_),
    .ZN(_11017_));
 AND4_X1 _16865_ (.A1(_10987_),
    .A2(_10996_),
    .A3(_11007_),
    .A4(_11017_),
    .ZN(_11018_));
 BUF_X4 _16866_ (.A(_11018_),
    .Z(_11019_));
 NOR4_X2 _16867_ (.A1(_10334_),
    .A2(_10374_),
    .A3(net18),
    .A4(_10923_),
    .ZN(_11020_));
 INV_X1 _16868_ (.A(_00139_),
    .ZN(_11021_));
 MUX2_X1 _16869_ (.A(_11021_),
    .B(_10451_),
    .S(_10386_),
    .Z(_11022_));
 AOI22_X1 _16870_ (.A1(_10976_),
    .A2(_11019_),
    .B1(_11020_),
    .B2(_11022_),
    .ZN(_11023_));
 OAI211_X2 _16871_ (.A(_10899_),
    .B(_10386_),
    .C1(_10387_),
    .C2(_10392_),
    .ZN(_11024_));
 AND2_X2 _16872_ (.A1(_11023_),
    .A2(_11024_),
    .ZN(_11025_));
 INV_X4 _16873_ (.A(_11025_),
    .ZN(_15864_));
 BUF_X8 _16874_ (.A(_11025_),
    .Z(_15860_));
 NOR2_X1 _16875_ (.A1(_10453_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .ZN(_11026_));
 AOI21_X1 _16876_ (.A(_11026_),
    .B1(_00310_),
    .B2(_10439_),
    .ZN(_11027_));
 INV_X1 _16877_ (.A(_00309_),
    .ZN(_11028_));
 AOI221_X2 _16878_ (.A(_10998_),
    .B1(_11027_),
    .B2(_10465_),
    .C1(_11028_),
    .C2(_10964_),
    .ZN(_11029_));
 MUX2_X1 _16879_ (.A(_00323_),
    .B(_00325_),
    .S(_10454_),
    .Z(_11030_));
 MUX2_X1 _16880_ (.A(_00324_),
    .B(_00326_),
    .S(_10454_),
    .Z(_11031_));
 MUX2_X1 _16881_ (.A(_11030_),
    .B(_11031_),
    .S(_10444_),
    .Z(_11032_));
 AOI21_X4 _16882_ (.A(_11029_),
    .B1(_11032_),
    .B2(_10995_),
    .ZN(_11033_));
 BUF_X4 _16883_ (.A(_10431_),
    .Z(_11034_));
 MUX2_X1 _16884_ (.A(_00315_),
    .B(_00319_),
    .S(_11034_),
    .Z(_11035_));
 MUX2_X1 _16885_ (.A(_00318_),
    .B(_00322_),
    .S(_11034_),
    .Z(_11036_));
 OAI22_X1 _16886_ (.A1(_10980_),
    .A2(_11035_),
    .B1(_11036_),
    .B2(_10977_),
    .ZN(_11037_));
 MUX2_X1 _16887_ (.A(_00316_),
    .B(_00320_),
    .S(_11034_),
    .Z(_11038_));
 MUX2_X1 _16888_ (.A(_00317_),
    .B(_00321_),
    .S(_11034_),
    .Z(_11039_));
 OAI22_X1 _16889_ (.A1(_10880_),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_10716_),
    .ZN(_11040_));
 OR3_X2 _16890_ (.A1(_10962_),
    .A2(_11037_),
    .A3(_11040_),
    .ZN(_11041_));
 NAND2_X2 _16891_ (.A1(_10451_),
    .A2(_10708_),
    .ZN(_11042_));
 MUX2_X1 _16892_ (.A(_00334_),
    .B(_00338_),
    .S(_11034_),
    .Z(_11043_));
 MUX2_X1 _16893_ (.A(_00332_),
    .B(_00336_),
    .S(_11034_),
    .Z(_11044_));
 OAI22_X1 _16894_ (.A1(_10977_),
    .A2(_11043_),
    .B1(_11044_),
    .B2(_10880_),
    .ZN(_11045_));
 MUX2_X1 _16895_ (.A(_00331_),
    .B(_00335_),
    .S(_11034_),
    .Z(_11046_));
 MUX2_X1 _16896_ (.A(_00333_),
    .B(_00337_),
    .S(_11034_),
    .Z(_11047_));
 OAI22_X1 _16897_ (.A1(_10980_),
    .A2(_11046_),
    .B1(_11047_),
    .B2(_10715_),
    .ZN(_11048_));
 OR3_X2 _16898_ (.A1(_11042_),
    .A2(_11045_),
    .A3(_11048_),
    .ZN(_11049_));
 MUX2_X1 _16899_ (.A(_00311_),
    .B(_00313_),
    .S(_10439_),
    .Z(_11050_));
 MUX2_X1 _16900_ (.A(_00312_),
    .B(_00314_),
    .S(_10439_),
    .Z(_11051_));
 MUX2_X1 _16901_ (.A(_11050_),
    .B(_11051_),
    .S(_10444_),
    .Z(_11052_));
 MUX2_X1 _16902_ (.A(_00327_),
    .B(_00329_),
    .S(_10457_),
    .Z(_11053_));
 MUX2_X1 _16903_ (.A(_00328_),
    .B(_00330_),
    .S(_10457_),
    .Z(_11054_));
 MUX2_X1 _16904_ (.A(_11053_),
    .B(_11054_),
    .S(_10465_),
    .Z(_11055_));
 AOI22_X4 _16905_ (.A1(_10988_),
    .A2(_11052_),
    .B1(_11055_),
    .B2(_11006_),
    .ZN(_11056_));
 NAND4_X4 _16906_ (.A1(_11033_),
    .A2(_11041_),
    .A3(_11049_),
    .A4(_11056_),
    .ZN(_11057_));
 MUX2_X1 _16907_ (.A(_00138_),
    .B(_10474_),
    .S(_10386_),
    .Z(_11058_));
 AND2_X2 _16908_ (.A1(_10326_),
    .A2(_10316_),
    .ZN(_11059_));
 NAND4_X4 _16909_ (.A1(_10389_),
    .A2(_10371_),
    .A3(_10375_),
    .A4(_11059_),
    .ZN(_11060_));
 OAI22_X4 _16910_ (.A1(_10974_),
    .A2(_11057_),
    .B1(_11058_),
    .B2(_11060_),
    .ZN(_11061_));
 INV_X1 _16911_ (.A(_10903_),
    .ZN(_11062_));
 AOI211_X2 _16912_ (.A(_11062_),
    .B(_10929_),
    .C1(_10930_),
    .C2(_10931_),
    .ZN(_11063_));
 NOR2_X2 _16913_ (.A1(_11061_),
    .A2(_11063_),
    .ZN(_11064_));
 INV_X4 _16914_ (.A(_11064_),
    .ZN(_15869_));
 BUF_X4 _16915_ (.A(_11064_),
    .Z(_11065_));
 BUF_X4 _16916_ (.A(_11065_),
    .Z(_15873_));
 NOR2_X1 _16917_ (.A1(_10920_),
    .A2(_15873_),
    .ZN(_15506_));
 BUF_X4 _16918_ (.A(_15515_),
    .Z(_11066_));
 NAND2_X4 _16919_ (.A1(_10972_),
    .A2(_10976_),
    .ZN(_11067_));
 MUX2_X1 _16920_ (.A(_10925_),
    .B(_10436_),
    .S(_10926_),
    .Z(_11068_));
 OAI221_X2 _16921_ (.A(_11059_),
    .B1(_11068_),
    .B2(_10334_),
    .C1(_10901_),
    .C2(_10393_),
    .ZN(_11069_));
 BUF_X4 _16922_ (.A(_11069_),
    .Z(_11070_));
 AOI21_X4 _16923_ (.A(_15864_),
    .B1(_11067_),
    .B2(_11070_),
    .ZN(_11071_));
 OAI21_X4 _16924_ (.A(_11066_),
    .B1(_10920_),
    .B2(_11071_),
    .ZN(_11072_));
 INV_X1 _16925_ (.A(_11072_),
    .ZN(_15507_));
 AOI21_X4 _16926_ (.A(_10373_),
    .B1(_10895_),
    .B2(_10368_),
    .ZN(_11073_));
 AOI22_X4 _16927_ (.A1(_10371_),
    .A2(_10375_),
    .B1(_10928_),
    .B2(_11073_),
    .ZN(_11074_));
 NAND2_X1 _16928_ (.A1(_10873_),
    .A2(_11059_),
    .ZN(_11075_));
 MUX2_X1 _16929_ (.A(_00353_),
    .B(_00355_),
    .S(_10406_),
    .Z(_11076_));
 MUX2_X1 _16930_ (.A(_00354_),
    .B(_00356_),
    .S(_10406_),
    .Z(_11077_));
 MUX2_X1 _16931_ (.A(_11076_),
    .B(_11077_),
    .S(_10414_),
    .Z(_11078_));
 AOI21_X1 _16932_ (.A(_10891_),
    .B1(_11078_),
    .B2(_10709_),
    .ZN(_11079_));
 NAND2_X1 _16933_ (.A1(_10454_),
    .A2(_00340_),
    .ZN(_11080_));
 OAI21_X1 _16934_ (.A(_11080_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .B2(net357),
    .ZN(_11081_));
 OAI22_X2 _16935_ (.A1(_00339_),
    .A2(_10716_),
    .B1(_11081_),
    .B2(_10696_),
    .ZN(_11082_));
 OAI21_X2 _16936_ (.A(_11079_),
    .B1(_11082_),
    .B2(_10709_),
    .ZN(_11083_));
 NAND3_X4 _16937_ (.A1(_11034_),
    .A2(_10421_),
    .A3(_10472_),
    .ZN(_11084_));
 MUX2_X1 _16938_ (.A(_00341_),
    .B(_00343_),
    .S(_10438_),
    .Z(_11085_));
 MUX2_X1 _16939_ (.A(_00342_),
    .B(_00344_),
    .S(_10438_),
    .Z(_11086_));
 MUX2_X1 _16940_ (.A(_11085_),
    .B(_11086_),
    .S(_10443_),
    .Z(_11087_));
 NOR2_X1 _16941_ (.A1(_11084_),
    .A2(_11087_),
    .ZN(_11088_));
 MUX2_X1 _16942_ (.A(_00345_),
    .B(_00349_),
    .S(_10984_),
    .Z(_11089_));
 MUX2_X1 _16943_ (.A(_00347_),
    .B(_00351_),
    .S(_10984_),
    .Z(_11090_));
 MUX2_X1 _16944_ (.A(_11089_),
    .B(_11090_),
    .S(_10439_),
    .Z(_11091_));
 NOR3_X1 _16945_ (.A1(_10444_),
    .A2(_10962_),
    .A3(_11091_),
    .ZN(_11092_));
 NOR2_X2 _16946_ (.A1(_11088_),
    .A2(_11092_),
    .ZN(_11093_));
 MUX2_X1 _16947_ (.A(_00362_),
    .B(_00366_),
    .S(_10431_),
    .Z(_11094_));
 MUX2_X1 _16948_ (.A(_00364_),
    .B(_00368_),
    .S(_10431_),
    .Z(_11095_));
 MUX2_X1 _16949_ (.A(_11094_),
    .B(_11095_),
    .S(_10454_),
    .Z(_11096_));
 NAND2_X4 _16950_ (.A1(_10443_),
    .A2(_10944_),
    .ZN(_11097_));
 NOR2_X1 _16951_ (.A1(_11096_),
    .A2(_11097_),
    .ZN(_11098_));
 NAND3_X4 _16952_ (.A1(_10431_),
    .A2(_10421_),
    .A3(_10872_),
    .ZN(_11099_));
 BUF_X4 _16953_ (.A(_10437_),
    .Z(_11100_));
 MUX2_X1 _16954_ (.A(_00357_),
    .B(_00359_),
    .S(_11100_),
    .Z(_11101_));
 MUX2_X1 _16955_ (.A(_00358_),
    .B(_00360_),
    .S(_11100_),
    .Z(_11102_));
 MUX2_X1 _16956_ (.A(_11101_),
    .B(_11102_),
    .S(_10443_),
    .Z(_11103_));
 NOR2_X1 _16957_ (.A1(_11099_),
    .A2(_11103_),
    .ZN(_11104_));
 NOR2_X2 _16958_ (.A1(_11098_),
    .A2(_11104_),
    .ZN(_11105_));
 MUX2_X1 _16959_ (.A(_00361_),
    .B(_00365_),
    .S(_10978_),
    .Z(_11106_));
 MUX2_X1 _16960_ (.A(_00363_),
    .B(_00367_),
    .S(_10978_),
    .Z(_11107_));
 MUX2_X1 _16961_ (.A(_11106_),
    .B(_11107_),
    .S(net401),
    .Z(_11108_));
 NOR3_X2 _16962_ (.A1(_10444_),
    .A2(_10473_),
    .A3(_11108_),
    .ZN(_11109_));
 MUX2_X1 _16963_ (.A(_00346_),
    .B(_00350_),
    .S(_10978_),
    .Z(_11110_));
 MUX2_X1 _16964_ (.A(_00348_),
    .B(_00352_),
    .S(_10978_),
    .Z(_11111_));
 MUX2_X1 _16965_ (.A(_11110_),
    .B(_11111_),
    .S(net401),
    .Z(_11112_));
 NOR3_X1 _16966_ (.A1(_10696_),
    .A2(_10709_),
    .A3(_11112_),
    .ZN(_11113_));
 OAI21_X2 _16967_ (.A(_10451_),
    .B1(_11109_),
    .B2(_11113_),
    .ZN(_11114_));
 AND4_X2 _16968_ (.A1(_11083_),
    .A2(_11093_),
    .A3(_11105_),
    .A4(_11114_),
    .ZN(_11115_));
 OAI22_X4 _16969_ (.A1(_11074_),
    .A2(_11075_),
    .B1(_11115_),
    .B2(_10974_),
    .ZN(_11116_));
 BUF_X4 _16970_ (.A(_11116_),
    .Z(_15876_));
 INV_X4 _16971_ (.A(_15876_),
    .ZN(_15880_));
 OR2_X1 _16972_ (.A1(_10412_),
    .A2(_10471_),
    .ZN(_11117_));
 MUX2_X1 _16973_ (.A(_00375_),
    .B(_00377_),
    .S(_10405_),
    .Z(_11118_));
 NOR2_X1 _16974_ (.A1(_11117_),
    .A2(_11118_),
    .ZN(_11119_));
 NAND2_X1 _16975_ (.A1(_10879_),
    .A2(_10707_),
    .ZN(_11120_));
 MUX2_X1 _16976_ (.A(_00392_),
    .B(_00394_),
    .S(_10456_),
    .Z(_11121_));
 OAI211_X2 _16977_ (.A(_10435_),
    .B(_10419_),
    .C1(_11120_),
    .C2(_11121_),
    .ZN(_11122_));
 MUX2_X1 _16978_ (.A(_00376_),
    .B(_00378_),
    .S(_10408_),
    .Z(_11123_));
 NOR3_X2 _16979_ (.A1(_10695_),
    .A2(_10872_),
    .A3(_11123_),
    .ZN(_11124_));
 MUX2_X1 _16980_ (.A(_00391_),
    .B(_00393_),
    .S(_10408_),
    .Z(_11125_));
 NOR3_X2 _16981_ (.A1(_10442_),
    .A2(_10472_),
    .A3(_11125_),
    .ZN(_11126_));
 NOR4_X4 _16982_ (.A1(_11119_),
    .A2(_11122_),
    .A3(_11124_),
    .A4(_11126_),
    .ZN(_11127_));
 MUX2_X1 _16983_ (.A(_00388_),
    .B(_00390_),
    .S(_10437_),
    .Z(_11128_));
 NOR2_X1 _16984_ (.A1(_11120_),
    .A2(_11128_),
    .ZN(_11129_));
 MUX2_X1 _16985_ (.A(_00387_),
    .B(_00389_),
    .S(_10404_),
    .Z(_11130_));
 NOR3_X2 _16986_ (.A1(_10879_),
    .A2(_10472_),
    .A3(_11130_),
    .ZN(_11131_));
 MUX2_X1 _16987_ (.A(_00372_),
    .B(_00374_),
    .S(_10404_),
    .Z(_11132_));
 NOR3_X2 _16988_ (.A1(_10694_),
    .A2(_10872_),
    .A3(_11132_),
    .ZN(_11133_));
 MUX2_X1 _16989_ (.A(_00371_),
    .B(_00373_),
    .S(_10404_),
    .Z(_11134_));
 OAI211_X2 _16990_ (.A(_10984_),
    .B(_10420_),
    .C1(_11117_),
    .C2(_11134_),
    .ZN(_11135_));
 NOR4_X4 _16991_ (.A1(_11129_),
    .A2(_11131_),
    .A3(_11133_),
    .A4(_11135_),
    .ZN(_11136_));
 MUX2_X1 _16992_ (.A(_00379_),
    .B(_00381_),
    .S(_10456_),
    .Z(_11137_));
 NOR2_X1 _16993_ (.A1(_10442_),
    .A2(_11137_),
    .ZN(_11138_));
 MUX2_X1 _16994_ (.A(_00380_),
    .B(_00382_),
    .S(_10408_),
    .Z(_11139_));
 NOR2_X1 _16995_ (.A1(_10695_),
    .A2(_11139_),
    .ZN(_11140_));
 NAND3_X1 _16996_ (.A1(_10431_),
    .A2(_10419_),
    .A3(_10472_),
    .ZN(_11141_));
 NAND2_X2 _16997_ (.A1(_10984_),
    .A2(_10944_),
    .ZN(_11142_));
 MUX2_X1 _16998_ (.A(_00395_),
    .B(_00397_),
    .S(_10404_),
    .Z(_11143_));
 NOR2_X1 _16999_ (.A1(_10879_),
    .A2(_11143_),
    .ZN(_11144_));
 MUX2_X1 _17000_ (.A(_00396_),
    .B(_00398_),
    .S(_10404_),
    .Z(_11145_));
 NOR2_X1 _17001_ (.A1(_10694_),
    .A2(_11145_),
    .ZN(_11146_));
 OAI33_X1 _17002_ (.A1(_11138_),
    .A2(_11140_),
    .A3(_11141_),
    .B1(_11142_),
    .B2(_11144_),
    .B3(_11146_),
    .ZN(_11147_));
 NAND2_X1 _17003_ (.A1(_10708_),
    .A2(_10997_),
    .ZN(_11148_));
 MUX2_X1 _17004_ (.A(_00383_),
    .B(_00385_),
    .S(_10408_),
    .Z(_11149_));
 NOR2_X1 _17005_ (.A1(_10879_),
    .A2(_11149_),
    .ZN(_11150_));
 MUX2_X1 _17006_ (.A(_00384_),
    .B(_00386_),
    .S(_10404_),
    .Z(_11151_));
 NOR2_X1 _17007_ (.A1(_10694_),
    .A2(_11151_),
    .ZN(_11152_));
 NOR3_X1 _17008_ (.A1(_10879_),
    .A2(_10336_),
    .A3(_00369_),
    .ZN(_11153_));
 NOR2_X1 _17009_ (.A1(_10456_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .ZN(_11154_));
 AND2_X1 _17010_ (.A1(_10408_),
    .A2(_00370_),
    .ZN(_11155_));
 NOR3_X1 _17011_ (.A1(_10694_),
    .A2(_11154_),
    .A3(_11155_),
    .ZN(_11156_));
 OAI33_X1 _17012_ (.A1(_11148_),
    .A2(_11150_),
    .A3(_11152_),
    .B1(_11153_),
    .B2(_11156_),
    .B3(_10998_),
    .ZN(_11157_));
 NOR4_X4 _17013_ (.A1(_11127_),
    .A2(_11136_),
    .A3(_11147_),
    .A4(_11157_),
    .ZN(_11158_));
 NAND2_X1 _17014_ (.A1(_10976_),
    .A2(_11158_),
    .ZN(_11159_));
 NAND3_X2 _17015_ (.A1(_10874_),
    .A2(_10386_),
    .A3(_11059_),
    .ZN(_11160_));
 NAND2_X1 _17016_ (.A1(_10326_),
    .A2(_10334_),
    .ZN(_11161_));
 AOI21_X4 _17017_ (.A(_11161_),
    .B1(_10375_),
    .B2(_10371_),
    .ZN(_11162_));
 OR2_X1 _17018_ (.A1(_10538_),
    .A2(_10386_),
    .ZN(_11163_));
 OAI221_X2 _17019_ (.A(_11159_),
    .B1(_11160_),
    .B2(_11162_),
    .C1(_11060_),
    .C2(_11163_),
    .ZN(_11164_));
 BUF_X4 _17020_ (.A(_11164_),
    .Z(_15884_));
 INV_X2 _17021_ (.A(_15884_),
    .ZN(_15888_));
 MUX2_X1 _17022_ (.A(_00413_),
    .B(_00415_),
    .S(_10710_),
    .Z(_11165_));
 NOR2_X1 _17023_ (.A1(_10444_),
    .A2(_11165_),
    .ZN(_11166_));
 MUX2_X1 _17024_ (.A(_00414_),
    .B(_00416_),
    .S(_10710_),
    .Z(_11167_));
 NOR2_X1 _17025_ (.A1(_10696_),
    .A2(_11167_),
    .ZN(_11168_));
 NOR3_X1 _17026_ (.A1(_10465_),
    .A2(_10337_),
    .A3(_00399_),
    .ZN(_11169_));
 NOR2_X1 _17027_ (.A1(_10439_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .ZN(_11170_));
 AND2_X1 _17028_ (.A1(_10710_),
    .A2(_00400_),
    .ZN(_11171_));
 NOR3_X1 _17029_ (.A1(_10696_),
    .A2(_11170_),
    .A3(_11171_),
    .ZN(_11172_));
 OAI33_X1 _17030_ (.A1(_11148_),
    .A2(_11166_),
    .A3(_11168_),
    .B1(_11169_),
    .B2(_11172_),
    .B3(_10998_),
    .ZN(_11173_));
 MUX2_X1 _17031_ (.A(_00406_),
    .B(_00410_),
    .S(_10431_),
    .Z(_11174_));
 NOR3_X2 _17032_ (.A1(_10696_),
    .A2(_10454_),
    .A3(_11174_),
    .ZN(_11175_));
 MUX2_X1 _17033_ (.A(_00408_),
    .B(_00412_),
    .S(_10431_),
    .Z(_11176_));
 MUX2_X1 _17034_ (.A(_00405_),
    .B(_00409_),
    .S(_10984_),
    .Z(_11177_));
 OAI22_X2 _17035_ (.A1(_10977_),
    .A2(_11176_),
    .B1(_11177_),
    .B2(_10980_),
    .ZN(_11178_));
 MUX2_X1 _17036_ (.A(_00407_),
    .B(_00411_),
    .S(_10984_),
    .Z(_11179_));
 NOR3_X2 _17037_ (.A1(_10414_),
    .A2(_10337_),
    .A3(_11179_),
    .ZN(_11180_));
 NOR4_X4 _17038_ (.A1(_10962_),
    .A2(_11175_),
    .A3(_11178_),
    .A4(_11180_),
    .ZN(_11181_));
 MUX2_X1 _17039_ (.A(_00418_),
    .B(_00420_),
    .S(_10406_),
    .Z(_11182_));
 NOR2_X1 _17040_ (.A1(_10696_),
    .A2(_11182_),
    .ZN(_11183_));
 MUX2_X1 _17041_ (.A(_00417_),
    .B(_00419_),
    .S(_10406_),
    .Z(_11184_));
 NOR2_X1 _17042_ (.A1(_10465_),
    .A2(_11184_),
    .ZN(_11185_));
 BUF_X4 _17043_ (.A(_10695_),
    .Z(_11186_));
 MUX2_X1 _17044_ (.A(_00402_),
    .B(_00404_),
    .S(_11100_),
    .Z(_11187_));
 NOR2_X1 _17045_ (.A1(_11186_),
    .A2(_11187_),
    .ZN(_11188_));
 MUX2_X1 _17046_ (.A(_00401_),
    .B(_00403_),
    .S(_11100_),
    .Z(_11189_));
 NOR2_X1 _17047_ (.A1(_10414_),
    .A2(_11189_),
    .ZN(_11190_));
 OAI33_X1 _17048_ (.A1(_11099_),
    .A2(_11183_),
    .A3(_11185_),
    .B1(_11188_),
    .B2(_11190_),
    .B3(_11084_),
    .ZN(_11191_));
 MUX2_X1 _17049_ (.A(_00425_),
    .B(_00427_),
    .S(_10438_),
    .Z(_11192_));
 NOR2_X1 _17050_ (.A1(_10465_),
    .A2(_11192_),
    .ZN(_11193_));
 MUX2_X1 _17051_ (.A(_00426_),
    .B(_00428_),
    .S(_10438_),
    .Z(_11194_));
 NOR2_X1 _17052_ (.A1(_11186_),
    .A2(_11194_),
    .ZN(_11195_));
 MUX2_X1 _17053_ (.A(_00421_),
    .B(_00423_),
    .S(_11100_),
    .Z(_11196_));
 NOR2_X1 _17054_ (.A1(_10414_),
    .A2(_11196_),
    .ZN(_11197_));
 MUX2_X1 _17055_ (.A(_00422_),
    .B(_00424_),
    .S(_10457_),
    .Z(_11198_));
 NOR2_X1 _17056_ (.A1(_11186_),
    .A2(_11198_),
    .ZN(_11199_));
 NAND2_X1 _17057_ (.A1(_10435_),
    .A2(_10944_),
    .ZN(_11200_));
 OAI33_X1 _17058_ (.A1(_11142_),
    .A2(_11193_),
    .A3(_11195_),
    .B1(_11197_),
    .B2(_11199_),
    .B3(_11200_),
    .ZN(_11201_));
 NOR4_X4 _17059_ (.A1(_11173_),
    .A2(_11201_),
    .A3(_11191_),
    .A4(_11181_),
    .ZN(_11202_));
 NAND2_X1 _17060_ (.A1(_10976_),
    .A2(_11202_),
    .ZN(_11203_));
 NAND2_X1 _17061_ (.A1(_10500_),
    .A2(_11059_),
    .ZN(_11204_));
 OAI21_X4 _17062_ (.A(_11203_),
    .B1(_11204_),
    .B2(_11074_),
    .ZN(_15892_));
 INV_X4 _17063_ (.A(_15892_),
    .ZN(_15896_));
 MUX2_X1 _17064_ (.A(_00452_),
    .B(_00456_),
    .S(_10430_),
    .Z(_11205_));
 MUX2_X1 _17065_ (.A(_00454_),
    .B(_00458_),
    .S(_10430_),
    .Z(_11206_));
 MUX2_X1 _17066_ (.A(_11205_),
    .B(_11206_),
    .S(_11100_),
    .Z(_11207_));
 MUX2_X1 _17067_ (.A(_00436_),
    .B(_00440_),
    .S(_10430_),
    .Z(_11208_));
 MUX2_X1 _17068_ (.A(_00438_),
    .B(_00442_),
    .S(_10430_),
    .Z(_11209_));
 MUX2_X1 _17069_ (.A(_11208_),
    .B(_11209_),
    .S(_11100_),
    .Z(_11210_));
 MUX2_X1 _17070_ (.A(_11207_),
    .B(_11210_),
    .S(_10473_),
    .Z(_11211_));
 MUX2_X1 _17071_ (.A(_00437_),
    .B(_00453_),
    .S(_10707_),
    .Z(_11212_));
 MUX2_X1 _17072_ (.A(_00441_),
    .B(_00457_),
    .S(_10707_),
    .Z(_11213_));
 MUX2_X1 _17073_ (.A(_11212_),
    .B(_11213_),
    .S(_10984_),
    .Z(_11214_));
 MUX2_X1 _17074_ (.A(_00435_),
    .B(_00451_),
    .S(_10707_),
    .Z(_11215_));
 MUX2_X1 _17075_ (.A(_00439_),
    .B(_00455_),
    .S(_10707_),
    .Z(_11216_));
 MUX2_X1 _17076_ (.A(_11215_),
    .B(_11216_),
    .S(_10431_),
    .Z(_11217_));
 MUX2_X1 _17077_ (.A(_11214_),
    .B(_11217_),
    .S(_10337_),
    .Z(_11218_));
 NAND2_X1 _17078_ (.A1(_10696_),
    .A2(_10451_),
    .ZN(_11219_));
 OAI22_X4 _17079_ (.A1(_11015_),
    .A2(_11211_),
    .B1(_11218_),
    .B2(_11219_),
    .ZN(_11220_));
 MUX2_X1 _17080_ (.A(_00443_),
    .B(_00445_),
    .S(_10409_),
    .Z(_11221_));
 NOR2_X1 _17081_ (.A1(_10941_),
    .A2(_11221_),
    .ZN(_11222_));
 MUX2_X1 _17082_ (.A(_00444_),
    .B(_00446_),
    .S(_10405_),
    .Z(_11223_));
 NOR2_X1 _17083_ (.A1(_11186_),
    .A2(_11223_),
    .ZN(_11224_));
 NOR3_X1 _17084_ (.A1(_10473_),
    .A2(_11222_),
    .A3(_11224_),
    .ZN(_11225_));
 INV_X1 _17085_ (.A(_00429_),
    .ZN(_11226_));
 NOR2_X1 _17086_ (.A1(_10437_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .ZN(_11227_));
 AOI21_X1 _17087_ (.A(_11227_),
    .B1(_00430_),
    .B2(net397),
    .ZN(_11228_));
 AOI221_X2 _17088_ (.A(_10708_),
    .B1(_11226_),
    .B2(_10964_),
    .C1(_11228_),
    .C2(_10442_),
    .ZN(_11229_));
 MUX2_X1 _17089_ (.A(_00447_),
    .B(_00449_),
    .S(_10405_),
    .Z(_11230_));
 NOR2_X1 _17090_ (.A1(_10941_),
    .A2(_11230_),
    .ZN(_11231_));
 MUX2_X1 _17091_ (.A(_00448_),
    .B(_00450_),
    .S(_10437_),
    .Z(_11232_));
 NOR2_X1 _17092_ (.A1(_10695_),
    .A2(_11232_),
    .ZN(_11233_));
 NOR3_X1 _17093_ (.A1(_10473_),
    .A2(_11231_),
    .A3(_11233_),
    .ZN(_11234_));
 MUX2_X1 _17094_ (.A(_00431_),
    .B(_00433_),
    .S(_10437_),
    .Z(_11235_));
 NOR2_X1 _17095_ (.A1(_10413_),
    .A2(_11235_),
    .ZN(_11236_));
 MUX2_X1 _17096_ (.A(_00432_),
    .B(_00434_),
    .S(_10437_),
    .Z(_11237_));
 NOR2_X1 _17097_ (.A1(_10695_),
    .A2(_11237_),
    .ZN(_11238_));
 NOR3_X1 _17098_ (.A1(_10708_),
    .A2(_11236_),
    .A3(_11238_),
    .ZN(_11239_));
 OAI33_X1 _17099_ (.A1(_10891_),
    .A2(_11225_),
    .A3(_11229_),
    .B1(_11234_),
    .B2(_11239_),
    .B3(_10881_),
    .ZN(_11240_));
 NOR2_X4 _17100_ (.A1(_11220_),
    .A2(_11240_),
    .ZN(_11241_));
 NOR2_X1 _17101_ (.A1(_10974_),
    .A2(_11241_),
    .ZN(_11242_));
 NOR2_X2 _17102_ (.A1(_10923_),
    .A2(_11074_),
    .ZN(_11243_));
 AOI21_X4 _17103_ (.A(_11242_),
    .B1(_11243_),
    .B2(_10501_),
    .ZN(_15904_));
 NAND2_X1 _17104_ (.A1(_10502_),
    .A2(_11243_),
    .ZN(_11244_));
 MUX2_X1 _17105_ (.A(_00465_),
    .B(_00481_),
    .S(_10872_),
    .Z(_11245_));
 MUX2_X1 _17106_ (.A(_00469_),
    .B(_00485_),
    .S(_10872_),
    .Z(_11246_));
 MUX2_X1 _17107_ (.A(_11245_),
    .B(_11246_),
    .S(_11034_),
    .Z(_11247_));
 NAND3_X4 _17108_ (.A1(_10696_),
    .A2(_10337_),
    .A3(_10451_),
    .ZN(_11248_));
 NAND3_X4 _17109_ (.A1(_11186_),
    .A2(_10454_),
    .A3(_10451_),
    .ZN(_11249_));
 MUX2_X1 _17110_ (.A(_00467_),
    .B(_00483_),
    .S(_10707_),
    .Z(_11250_));
 MUX2_X1 _17111_ (.A(_00471_),
    .B(_00487_),
    .S(_10707_),
    .Z(_11251_));
 MUX2_X1 _17112_ (.A(_11250_),
    .B(_11251_),
    .S(_10685_),
    .Z(_11252_));
 OAI22_X4 _17113_ (.A1(_11247_),
    .A2(_11248_),
    .B1(_11249_),
    .B2(_11252_),
    .ZN(_11253_));
 MUX2_X1 _17114_ (.A(_00477_),
    .B(_00479_),
    .S(_10409_),
    .Z(_11254_));
 MUX2_X1 _17115_ (.A(_00478_),
    .B(_00480_),
    .S(_10409_),
    .Z(_11255_));
 MUX2_X1 _17116_ (.A(_11254_),
    .B(_11255_),
    .S(_10413_),
    .Z(_11256_));
 MUX2_X1 _17117_ (.A(_00461_),
    .B(_00463_),
    .S(_10405_),
    .Z(_11257_));
 MUX2_X1 _17118_ (.A(_00462_),
    .B(_00464_),
    .S(_10405_),
    .Z(_11258_));
 MUX2_X1 _17119_ (.A(_11257_),
    .B(_11258_),
    .S(_10413_),
    .Z(_11259_));
 OAI22_X4 _17120_ (.A1(_11099_),
    .A2(_11256_),
    .B1(_11259_),
    .B2(_11084_),
    .ZN(_11260_));
 MUX2_X1 _17121_ (.A(_00482_),
    .B(_00486_),
    .S(_10684_),
    .Z(_11261_));
 MUX2_X1 _17122_ (.A(_00484_),
    .B(_00488_),
    .S(_10684_),
    .Z(_11262_));
 MUX2_X1 _17123_ (.A(_11261_),
    .B(_11262_),
    .S(_10710_),
    .Z(_11263_));
 MUX2_X1 _17124_ (.A(_00466_),
    .B(_00470_),
    .S(_10434_),
    .Z(_11264_));
 MUX2_X1 _17125_ (.A(_00468_),
    .B(_00472_),
    .S(_10434_),
    .Z(_11265_));
 MUX2_X1 _17126_ (.A(_11264_),
    .B(_11265_),
    .S(_10453_),
    .Z(_11266_));
 NOR2_X2 _17127_ (.A1(_10421_),
    .A2(_10708_),
    .ZN(_11267_));
 NAND2_X2 _17128_ (.A1(_10443_),
    .A2(_11267_),
    .ZN(_11268_));
 OAI22_X4 _17129_ (.A1(_11097_),
    .A2(_11263_),
    .B1(_11266_),
    .B2(_11268_),
    .ZN(_11269_));
 NOR2_X1 _17130_ (.A1(net334),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .ZN(_11270_));
 AOI21_X1 _17131_ (.A(_11270_),
    .B1(_00460_),
    .B2(_10409_),
    .ZN(_11271_));
 NAND2_X1 _17132_ (.A1(_10442_),
    .A2(_11271_),
    .ZN(_11272_));
 INV_X1 _17133_ (.A(_00459_),
    .ZN(_11273_));
 AOI21_X1 _17134_ (.A(_10707_),
    .B1(_11273_),
    .B2(_10964_),
    .ZN(_11274_));
 MUX2_X1 _17135_ (.A(_00473_),
    .B(_00475_),
    .S(_10404_),
    .Z(_11275_));
 MUX2_X1 _17136_ (.A(_00474_),
    .B(_00476_),
    .S(_10404_),
    .Z(_11276_));
 MUX2_X1 _17137_ (.A(_11275_),
    .B(_11276_),
    .S(_10412_),
    .Z(_11277_));
 AOI221_X2 _17138_ (.A(_10891_),
    .B1(_11272_),
    .B2(_11274_),
    .C1(_11277_),
    .C2(_10708_),
    .ZN(_11278_));
 NOR4_X4 _17139_ (.A1(_11253_),
    .A2(_11260_),
    .A3(_11269_),
    .A4(_11278_),
    .ZN(_11279_));
 OAI21_X4 _17140_ (.A(_11244_),
    .B1(_11279_),
    .B2(_10974_),
    .ZN(_15908_));
 INV_X1 _17141_ (.A(_15908_),
    .ZN(_15912_));
 NOR2_X1 _17142_ (.A1(_10452_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .ZN(_11280_));
 AOI21_X1 _17143_ (.A(_11280_),
    .B1(_00490_),
    .B2(_10438_),
    .ZN(_11281_));
 INV_X1 _17144_ (.A(_00489_),
    .ZN(_11282_));
 AOI221_X2 _17145_ (.A(_10998_),
    .B1(_11281_),
    .B2(_10413_),
    .C1(_11282_),
    .C2(_10964_),
    .ZN(_11283_));
 MUX2_X1 _17146_ (.A(_00503_),
    .B(_00505_),
    .S(_10438_),
    .Z(_11284_));
 MUX2_X1 _17147_ (.A(_00504_),
    .B(_00506_),
    .S(_10438_),
    .Z(_11285_));
 MUX2_X1 _17148_ (.A(_11284_),
    .B(_11285_),
    .S(_10443_),
    .Z(_11286_));
 MUX2_X1 _17149_ (.A(_00495_),
    .B(_00499_),
    .S(_10685_),
    .Z(_11287_));
 NOR2_X1 _17150_ (.A1(_10980_),
    .A2(_11287_),
    .ZN(_11288_));
 MUX2_X1 _17151_ (.A(_00496_),
    .B(_00500_),
    .S(_10984_),
    .Z(_11289_));
 NOR3_X1 _17152_ (.A1(_11186_),
    .A2(_10439_),
    .A3(_11289_),
    .ZN(_11290_));
 MUX2_X1 _17153_ (.A(_00498_),
    .B(_00502_),
    .S(_10984_),
    .Z(_11291_));
 NOR2_X1 _17154_ (.A1(_10977_),
    .A2(_11291_),
    .ZN(_11292_));
 MUX2_X1 _17155_ (.A(_00497_),
    .B(_00501_),
    .S(_10978_),
    .Z(_11293_));
 NOR3_X1 _17156_ (.A1(_10443_),
    .A2(_10337_),
    .A3(_11293_),
    .ZN(_11294_));
 NOR4_X2 _17157_ (.A1(_11288_),
    .A2(_11290_),
    .A3(_11292_),
    .A4(_11294_),
    .ZN(_11295_));
 AOI221_X2 _17158_ (.A(_11283_),
    .B1(_11286_),
    .B2(_10995_),
    .C1(_11295_),
    .C2(_11267_),
    .ZN(_11296_));
 MUX2_X1 _17159_ (.A(_00515_),
    .B(_00517_),
    .S(_11100_),
    .Z(_11297_));
 NOR2_X1 _17160_ (.A1(_10443_),
    .A2(_11297_),
    .ZN(_11298_));
 MUX2_X1 _17161_ (.A(_00516_),
    .B(_00518_),
    .S(net397),
    .Z(_11299_));
 NOR2_X1 _17162_ (.A1(_11186_),
    .A2(_11299_),
    .ZN(_11300_));
 MUX2_X1 _17163_ (.A(_00511_),
    .B(_00513_),
    .S(net397),
    .Z(_11301_));
 NOR2_X1 _17164_ (.A1(_10941_),
    .A2(_11301_),
    .ZN(_11302_));
 MUX2_X1 _17165_ (.A(_00512_),
    .B(_00514_),
    .S(_10409_),
    .Z(_11303_));
 NOR2_X1 _17166_ (.A1(_11186_),
    .A2(_11303_),
    .ZN(_11304_));
 OAI33_X1 _17167_ (.A1(_11142_),
    .A2(_11298_),
    .A3(_11300_),
    .B1(_11302_),
    .B2(_11304_),
    .B3(_11200_),
    .ZN(_11305_));
 MUX2_X1 _17168_ (.A(_00507_),
    .B(_00509_),
    .S(_11100_),
    .Z(_11306_));
 MUX2_X1 _17169_ (.A(_00508_),
    .B(_00510_),
    .S(_11100_),
    .Z(_11307_));
 MUX2_X1 _17170_ (.A(_11306_),
    .B(_11307_),
    .S(_10443_),
    .Z(_11308_));
 MUX2_X1 _17171_ (.A(_00491_),
    .B(_00493_),
    .S(_10453_),
    .Z(_11309_));
 MUX2_X1 _17172_ (.A(_00492_),
    .B(_00494_),
    .S(_10453_),
    .Z(_11310_));
 MUX2_X1 _17173_ (.A(_11309_),
    .B(_11310_),
    .S(_10465_),
    .Z(_11311_));
 AOI221_X2 _17174_ (.A(_11305_),
    .B1(_11308_),
    .B2(_11006_),
    .C1(_11311_),
    .C2(_10988_),
    .ZN(_11312_));
 NAND2_X4 _17175_ (.A1(_11296_),
    .A2(_11312_),
    .ZN(_11313_));
 NAND2_X1 _17176_ (.A1(_10498_),
    .A2(_11059_),
    .ZN(_11314_));
 OAI22_X4 _17177_ (.A1(_10974_),
    .A2(_11313_),
    .B1(_11314_),
    .B2(_11074_),
    .ZN(_15916_));
 INV_X4 _17178_ (.A(_15916_),
    .ZN(_15920_));
 INV_X4 _17179_ (.A(_10902_),
    .ZN(_11315_));
 AOI21_X1 _17180_ (.A(_10509_),
    .B1(_10330_),
    .B2(_10385_),
    .ZN(_11316_));
 NAND2_X1 _17181_ (.A1(_00140_),
    .A2(_10330_),
    .ZN(_11317_));
 OAI21_X1 _17182_ (.A(_11073_),
    .B1(_10353_),
    .B2(_11317_),
    .ZN(_11318_));
 OAI22_X2 _17183_ (.A1(_11315_),
    .A2(_11073_),
    .B1(_11316_),
    .B2(_11318_),
    .ZN(_11319_));
 AOI211_X2 _17184_ (.A(_00174_),
    .B(_10334_),
    .C1(_10371_),
    .C2(_10375_),
    .ZN(_11320_));
 AOI221_X2 _17185_ (.A(_10403_),
    .B1(_10926_),
    .B2(_11319_),
    .C1(_11320_),
    .C2(_10928_),
    .ZN(_11321_));
 MUX2_X1 _17186_ (.A(_00527_),
    .B(_00543_),
    .S(_10872_),
    .Z(_11322_));
 MUX2_X1 _17187_ (.A(_00531_),
    .B(_00547_),
    .S(_10872_),
    .Z(_11323_));
 MUX2_X1 _17188_ (.A(_11322_),
    .B(_11323_),
    .S(_10432_),
    .Z(_11324_));
 MUX2_X1 _17189_ (.A(_00525_),
    .B(_00541_),
    .S(_10872_),
    .Z(_11325_));
 MUX2_X1 _17190_ (.A(_00529_),
    .B(_00545_),
    .S(_10872_),
    .Z(_11326_));
 MUX2_X1 _17191_ (.A(_11325_),
    .B(_11326_),
    .S(_10432_),
    .Z(_11327_));
 OAI22_X4 _17192_ (.A1(_11249_),
    .A2(_11324_),
    .B1(_11327_),
    .B2(_11248_),
    .ZN(_11328_));
 MUX2_X1 _17193_ (.A(_00537_),
    .B(_00539_),
    .S(net397),
    .Z(_11329_));
 MUX2_X1 _17194_ (.A(_00538_),
    .B(_00540_),
    .S(net397),
    .Z(_11330_));
 MUX2_X1 _17195_ (.A(_11329_),
    .B(_11330_),
    .S(_10941_),
    .Z(_11331_));
 MUX2_X1 _17196_ (.A(_00521_),
    .B(_00523_),
    .S(net401),
    .Z(_11332_));
 MUX2_X1 _17197_ (.A(_00522_),
    .B(_00524_),
    .S(net401),
    .Z(_11333_));
 MUX2_X1 _17198_ (.A(_11332_),
    .B(_11333_),
    .S(_10941_),
    .Z(_11334_));
 OAI22_X4 _17199_ (.A1(_11099_),
    .A2(_11331_),
    .B1(_11334_),
    .B2(_11084_),
    .ZN(_11335_));
 MUX2_X1 _17200_ (.A(_00542_),
    .B(_00546_),
    .S(_10978_),
    .Z(_11336_));
 MUX2_X1 _17201_ (.A(_00544_),
    .B(_00548_),
    .S(_10978_),
    .Z(_11337_));
 MUX2_X1 _17202_ (.A(_11336_),
    .B(_11337_),
    .S(net397),
    .Z(_11338_));
 MUX2_X1 _17203_ (.A(_00526_),
    .B(_00530_),
    .S(_10684_),
    .Z(_11339_));
 MUX2_X1 _17204_ (.A(_00528_),
    .B(_00532_),
    .S(_10978_),
    .Z(_11340_));
 MUX2_X1 _17205_ (.A(_11339_),
    .B(_11340_),
    .S(net397),
    .Z(_11341_));
 OAI22_X4 _17206_ (.A1(_11097_),
    .A2(_11338_),
    .B1(_11341_),
    .B2(_11268_),
    .ZN(_11342_));
 NAND2_X1 _17207_ (.A1(_10453_),
    .A2(_00520_),
    .ZN(_11343_));
 OAI21_X1 _17208_ (.A(_11343_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B2(net397),
    .ZN(_11344_));
 OAI221_X1 _17209_ (.A(_10473_),
    .B1(_00519_),
    .B2(_10715_),
    .C1(_11344_),
    .C2(_11186_),
    .ZN(_11345_));
 MUX2_X1 _17210_ (.A(_00533_),
    .B(_00535_),
    .S(net334),
    .Z(_11346_));
 MUX2_X1 _17211_ (.A(_00534_),
    .B(_00536_),
    .S(net334),
    .Z(_11347_));
 MUX2_X1 _17212_ (.A(_11346_),
    .B(_11347_),
    .S(_10879_),
    .Z(_11348_));
 AOI21_X1 _17213_ (.A(_10891_),
    .B1(_11348_),
    .B2(_10709_),
    .ZN(_11349_));
 AND2_X2 _17214_ (.A1(_11345_),
    .A2(_11349_),
    .ZN(_11350_));
 OR4_X4 _17215_ (.A1(_11328_),
    .A2(_11335_),
    .A3(_11342_),
    .A4(_11350_),
    .ZN(_11351_));
 OAI21_X4 _17216_ (.A(_10673_),
    .B1(_10317_),
    .B2(_11351_),
    .ZN(_11352_));
 OR2_X1 _17217_ (.A1(_11321_),
    .A2(_11352_),
    .ZN(_11353_));
 BUF_X4 _17218_ (.A(_11353_),
    .Z(_15929_));
 INV_X2 _17219_ (.A(_15929_),
    .ZN(_15925_));
 INV_X2 _17220_ (.A(_15936_),
    .ZN(_15932_));
 OR2_X1 _17221_ (.A1(_10380_),
    .A2(_10898_),
    .ZN(_11354_));
 NAND3_X2 _17222_ (.A1(_10477_),
    .A2(_10661_),
    .A3(_11354_),
    .ZN(_15522_));
 INV_X1 _17223_ (.A(_15522_),
    .ZN(_15529_));
 NAND3_X4 _17224_ (.A1(_10488_),
    .A2(_10661_),
    .A3(_10898_),
    .ZN(_11355_));
 CLKBUF_X2 _17225_ (.A(_11355_),
    .Z(_11356_));
 BUF_X2 _17226_ (.A(_11356_),
    .Z(_15526_));
 BUF_X4 _17227_ (.A(_10567_),
    .Z(_11357_));
 BUF_X4 _17228_ (.A(_11357_),
    .Z(_11358_));
 NAND2_X1 _17229_ (.A1(_10621_),
    .A2(_00520_),
    .ZN(_11359_));
 OAI21_X1 _17230_ (.A(_11359_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B2(_10615_),
    .ZN(_11360_));
 OAI221_X1 _17231_ (.A(_11358_),
    .B1(_00519_),
    .B2(_10757_),
    .C1(_11360_),
    .C2(_10580_),
    .ZN(_11361_));
 BUF_X4 _17232_ (.A(_10790_),
    .Z(_11362_));
 BUF_X4 _17233_ (.A(_11362_),
    .Z(_11363_));
 MUX2_X1 _17234_ (.A(_00525_),
    .B(_00527_),
    .S(_11363_),
    .Z(_11364_));
 MUX2_X1 _17235_ (.A(_00526_),
    .B(_00528_),
    .S(_11363_),
    .Z(_11365_));
 BUF_X8 _17236_ (.A(_10862_),
    .Z(_11366_));
 MUX2_X1 _17237_ (.A(_11364_),
    .B(_11365_),
    .S(_11366_),
    .Z(_11367_));
 AOI21_X1 _17238_ (.A(_10830_),
    .B1(_11367_),
    .B2(_10766_),
    .ZN(_11368_));
 NAND2_X1 _17239_ (.A1(_11361_),
    .A2(_11368_),
    .ZN(_11369_));
 BUF_X8 _17240_ (.A(_10572_),
    .Z(_11370_));
 NAND2_X4 _17241_ (.A1(_10608_),
    .A2(_11370_),
    .ZN(_11371_));
 BUF_X8 _17242_ (.A(_10598_),
    .Z(_11372_));
 MUX2_X1 _17243_ (.A(_00541_),
    .B(_00543_),
    .S(_11372_),
    .Z(_11373_));
 MUX2_X1 _17244_ (.A(_00542_),
    .B(_00544_),
    .S(_11372_),
    .Z(_11374_));
 BUF_X4 _17245_ (.A(_10593_),
    .Z(_11375_));
 MUX2_X1 _17246_ (.A(_11373_),
    .B(_11374_),
    .S(_11375_),
    .Z(_11376_));
 MUX2_X1 _17247_ (.A(_00533_),
    .B(_00535_),
    .S(_11372_),
    .Z(_11377_));
 MUX2_X1 _17248_ (.A(_00534_),
    .B(_00536_),
    .S(_11372_),
    .Z(_11378_));
 MUX2_X1 _17249_ (.A(_11377_),
    .B(_11378_),
    .S(_11375_),
    .Z(_11379_));
 MUX2_X1 _17250_ (.A(_11376_),
    .B(_11379_),
    .S(_10569_),
    .Z(_11380_));
 MUX2_X1 _17251_ (.A(_00545_),
    .B(_00547_),
    .S(_10598_),
    .Z(_11381_));
 MUX2_X1 _17252_ (.A(_00546_),
    .B(_00548_),
    .S(_10598_),
    .Z(_11382_));
 BUF_X4 _17253_ (.A(_10592_),
    .Z(_11383_));
 MUX2_X1 _17254_ (.A(_11381_),
    .B(_11382_),
    .S(_11383_),
    .Z(_11384_));
 BUF_X4 _17255_ (.A(_10584_),
    .Z(_11385_));
 MUX2_X1 _17256_ (.A(_00537_),
    .B(_00539_),
    .S(_11385_),
    .Z(_11386_));
 MUX2_X1 _17257_ (.A(_00538_),
    .B(_00540_),
    .S(_11385_),
    .Z(_11387_));
 MUX2_X1 _17258_ (.A(_11386_),
    .B(_11387_),
    .S(_11383_),
    .Z(_11388_));
 MUX2_X1 _17259_ (.A(_11384_),
    .B(_11388_),
    .S(_10568_),
    .Z(_11389_));
 MUX2_X1 _17260_ (.A(_00529_),
    .B(_00531_),
    .S(_11385_),
    .Z(_11390_));
 MUX2_X1 _17261_ (.A(_00530_),
    .B(_00532_),
    .S(_11385_),
    .Z(_11391_));
 MUX2_X1 _17262_ (.A(_11390_),
    .B(_11391_),
    .S(_11383_),
    .Z(_11392_));
 MUX2_X1 _17263_ (.A(_00521_),
    .B(_00523_),
    .S(_11385_),
    .Z(_11393_));
 MUX2_X1 _17264_ (.A(_00522_),
    .B(_00524_),
    .S(_11385_),
    .Z(_11394_));
 MUX2_X1 _17265_ (.A(_11393_),
    .B(_11394_),
    .S(_11383_),
    .Z(_11395_));
 MUX2_X1 _17266_ (.A(_11392_),
    .B(_11395_),
    .S(_10568_),
    .Z(_11396_));
 MUX2_X1 _17267_ (.A(_11389_),
    .B(_11396_),
    .S(_10574_),
    .Z(_11397_));
 OAI221_X2 _17268_ (.A(_11369_),
    .B1(_11380_),
    .B2(_11371_),
    .C1(_11397_),
    .C2(_10609_),
    .ZN(_11398_));
 AND2_X1 _17269_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_10563_),
    .ZN(_11399_));
 AOI222_X2 _17270_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(_10741_),
    .B1(_10816_),
    .B2(_11398_),
    .C1(_11399_),
    .C2(_10870_),
    .ZN(_15928_));
 BUF_X1 _17271_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Z(_11400_));
 NOR3_X4 _17272_ (.A1(_10508_),
    .A2(_10912_),
    .A3(_10541_),
    .ZN(_11401_));
 OAI21_X4 _17273_ (.A(_11401_),
    .B1(_10677_),
    .B2(_10310_),
    .ZN(_11402_));
 NAND2_X1 _17274_ (.A1(_11400_),
    .A2(_11402_),
    .ZN(_11403_));
 NAND2_X1 _17275_ (.A1(_00555_),
    .A2(_11403_),
    .ZN(_11404_));
 NAND3_X2 _17276_ (.A1(_10873_),
    .A2(_10514_),
    .A3(_10917_),
    .ZN(_11405_));
 BUF_X4 _17277_ (.A(_11405_),
    .Z(_11406_));
 BUF_X4 _17278_ (.A(_11406_),
    .Z(_11407_));
 BUF_X4 _17279_ (.A(_11407_),
    .Z(_11408_));
 BUF_X4 _17280_ (.A(_11408_),
    .Z(_11409_));
 OR4_X1 _17281_ (.A1(_10373_),
    .A2(_10530_),
    .A3(_10531_),
    .A4(_10532_),
    .ZN(_11410_));
 NAND4_X1 _17282_ (.A1(_10508_),
    .A2(_10499_),
    .A3(_00174_),
    .A4(net284),
    .ZN(_11411_));
 NAND4_X1 _17283_ (.A1(_10508_),
    .A2(_00174_),
    .A3(_10538_),
    .A4(net283),
    .ZN(_11412_));
 AOI22_X2 _17284_ (.A1(_10522_),
    .A2(_11411_),
    .B1(_11412_),
    .B2(_10310_),
    .ZN(_11413_));
 OR3_X1 _17285_ (.A1(_10480_),
    .A2(_10549_),
    .A3(_10481_),
    .ZN(_11414_));
 AOI21_X1 _17286_ (.A(_10341_),
    .B1(_10522_),
    .B2(_10670_),
    .ZN(_11415_));
 AOI22_X2 _17287_ (.A1(_10342_),
    .A2(_10536_),
    .B1(_11415_),
    .B2(_10352_),
    .ZN(_11416_));
 OAI222_X2 _17288_ (.A1(_11410_),
    .A2(_10661_),
    .B1(_11413_),
    .B2(_11414_),
    .C1(_11416_),
    .C2(_10340_),
    .ZN(_11417_));
 NOR4_X4 _17289_ (.A1(_10894_),
    .A2(_10910_),
    .A3(_10918_),
    .A4(_11417_),
    .ZN(_11418_));
 CLKBUF_X3 _17290_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Z(_11419_));
 BUF_X4 _17291_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Z(_11420_));
 BUF_X4 _17292_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Z(_11421_));
 BUF_X4 _17293_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Z(_11422_));
 CLKBUF_X3 _17294_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_11423_));
 INV_X8 _17295_ (.A(_11423_),
    .ZN(_11424_));
 NOR3_X4 _17296_ (.A1(_11421_),
    .A2(_11422_),
    .A3(_11424_),
    .ZN(_11425_));
 NAND2_X4 _17297_ (.A1(_11420_),
    .A2(_11425_),
    .ZN(_11426_));
 NOR3_X4 _17298_ (.A1(_10305_),
    .A2(_11419_),
    .A3(_11426_),
    .ZN(_11427_));
 NAND2_X4 _17299_ (.A1(_11418_),
    .A2(_11427_),
    .ZN(_11428_));
 NOR3_X4 _17300_ (.A1(_10495_),
    .A2(_11409_),
    .A3(_11428_),
    .ZN(_11429_));
 MUX2_X1 _17301_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(_11404_),
    .S(_11429_),
    .Z(_00000_));
 BUF_X4 _17302_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(_11430_));
 BUF_X4 _17303_ (.A(_11400_),
    .Z(_11431_));
 BUF_X4 _17304_ (.A(_10402_),
    .Z(_11432_));
 AOI21_X4 _17305_ (.A(_11406_),
    .B1(_10670_),
    .B2(_11432_),
    .ZN(_11433_));
 AND2_X2 _17306_ (.A1(_11431_),
    .A2(_11433_),
    .ZN(_11434_));
 MUX2_X1 _17307_ (.A(_11430_),
    .B(_11434_),
    .S(_11429_),
    .Z(_00001_));
 INV_X1 _17308_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .ZN(_11435_));
 OAI22_X1 _17309_ (.A1(_11435_),
    .A2(_10565_),
    .B1(_10681_),
    .B2(_10397_),
    .ZN(_11436_));
 INV_X2 _17310_ (.A(_10792_),
    .ZN(_11437_));
 MUX2_X1 _17311_ (.A(_00262_),
    .B(_00264_),
    .S(_10621_),
    .Z(_11438_));
 MUX2_X1 _17312_ (.A(_00263_),
    .B(_00265_),
    .S(_10621_),
    .Z(_11439_));
 MUX2_X1 _17313_ (.A(_11438_),
    .B(_11439_),
    .S(_10629_),
    .Z(_11440_));
 AOI21_X1 _17314_ (.A(_11437_),
    .B1(_11440_),
    .B2(_10749_),
    .ZN(_11441_));
 NAND2_X1 _17315_ (.A1(_10616_),
    .A2(_00249_),
    .ZN(_11442_));
 OAI21_X1 _17316_ (.A(_11442_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .B2(_10616_),
    .ZN(_11443_));
 OAI22_X1 _17317_ (.A1(_00248_),
    .A2(_10758_),
    .B1(_11443_),
    .B2(_10582_),
    .ZN(_11444_));
 OAI21_X1 _17318_ (.A(_11441_),
    .B1(_11444_),
    .B2(_10750_),
    .ZN(_11445_));
 MUX2_X1 _17319_ (.A(_00270_),
    .B(_00272_),
    .S(_10614_),
    .Z(_11446_));
 MUX2_X1 _17320_ (.A(_00271_),
    .B(_00273_),
    .S(_10614_),
    .Z(_11447_));
 MUX2_X1 _17321_ (.A(_11446_),
    .B(_11447_),
    .S(_10797_),
    .Z(_11448_));
 MUX2_X1 _17322_ (.A(_00254_),
    .B(_00256_),
    .S(_10614_),
    .Z(_11449_));
 MUX2_X1 _17323_ (.A(_00255_),
    .B(_00257_),
    .S(_10614_),
    .Z(_11450_));
 MUX2_X1 _17324_ (.A(_11449_),
    .B(_11450_),
    .S(_10596_),
    .Z(_11451_));
 MUX2_X1 _17325_ (.A(_11448_),
    .B(_11451_),
    .S(_10576_),
    .Z(_11452_));
 NAND2_X4 _17326_ (.A1(_10608_),
    .A2(_10766_),
    .ZN(_11453_));
 BUF_X4 _17327_ (.A(_10858_),
    .Z(_11454_));
 MUX2_X1 _17328_ (.A(_00274_),
    .B(_00276_),
    .S(_11454_),
    .Z(_11455_));
 MUX2_X1 _17329_ (.A(_00275_),
    .B(_00277_),
    .S(_11454_),
    .Z(_11456_));
 MUX2_X1 _17330_ (.A(_11455_),
    .B(_11456_),
    .S(_11366_),
    .Z(_11457_));
 MUX2_X1 _17331_ (.A(_00258_),
    .B(_00260_),
    .S(_11454_),
    .Z(_11458_));
 MUX2_X1 _17332_ (.A(_00259_),
    .B(_00261_),
    .S(_11454_),
    .Z(_11459_));
 MUX2_X1 _17333_ (.A(_11458_),
    .B(_11459_),
    .S(_11366_),
    .Z(_11460_));
 MUX2_X1 _17334_ (.A(_11457_),
    .B(_11460_),
    .S(_10575_),
    .Z(_11461_));
 MUX2_X1 _17335_ (.A(_00266_),
    .B(_00268_),
    .S(_11454_),
    .Z(_11462_));
 MUX2_X1 _17336_ (.A(_00267_),
    .B(_00269_),
    .S(_11454_),
    .Z(_11463_));
 MUX2_X1 _17337_ (.A(_11462_),
    .B(_11463_),
    .S(_10595_),
    .Z(_11464_));
 MUX2_X1 _17338_ (.A(_00250_),
    .B(_00252_),
    .S(_11454_),
    .Z(_11465_));
 MUX2_X1 _17339_ (.A(_00251_),
    .B(_00253_),
    .S(_11454_),
    .Z(_11466_));
 MUX2_X1 _17340_ (.A(_11465_),
    .B(_11466_),
    .S(_10595_),
    .Z(_11467_));
 MUX2_X1 _17341_ (.A(_11464_),
    .B(_11467_),
    .S(_10575_),
    .Z(_11468_));
 MUX2_X1 _17342_ (.A(_11461_),
    .B(_11468_),
    .S(_10571_),
    .Z(_11469_));
 OAI221_X2 _17343_ (.A(_11445_),
    .B1(_11452_),
    .B2(_11453_),
    .C1(_10610_),
    .C2(_11469_),
    .ZN(_11470_));
 AOI21_X2 _17344_ (.A(_11436_),
    .B1(net293),
    .B2(_10565_),
    .ZN(_11471_));
 NOR3_X1 _17345_ (.A1(_00182_),
    .A2(_10565_),
    .A3(_10744_),
    .ZN(_11472_));
 AND2_X1 _17346_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_10565_),
    .ZN(_11473_));
 NOR3_X2 _17347_ (.A1(_10747_),
    .A2(_11472_),
    .A3(_11473_),
    .ZN(_11474_));
 NOR2_X4 _17348_ (.A1(_11471_),
    .A2(_11474_),
    .ZN(_15852_));
 INV_X2 _17349_ (.A(_15852_),
    .ZN(_15856_));
 BUF_X1 rebuffer21 (.A(_13061_),
    .Z(net292));
 INV_X2 _17351_ (.A(_15365_),
    .ZN(_11476_));
 OAI21_X1 _17352_ (.A(_10538_),
    .B1(_10499_),
    .B2(net315),
    .ZN(_11477_));
 NOR4_X2 _17353_ (.A1(_10549_),
    .A2(_10512_),
    .A3(_10912_),
    .A4(_11477_),
    .ZN(_11478_));
 NOR2_X1 _17354_ (.A1(_10480_),
    .A2(_10382_),
    .ZN(_11479_));
 OAI33_X1 _17355_ (.A1(_10305_),
    .A2(_10306_),
    .A3(_10384_),
    .B1(_10481_),
    .B2(_10484_),
    .B3(_10486_),
    .ZN(_11480_));
 AOI221_X2 _17356_ (.A(_11478_),
    .B1(_11479_),
    .B2(_11480_),
    .C1(_10487_),
    .C2(_10505_),
    .ZN(_11481_));
 BUF_X4 _17357_ (.A(_11481_),
    .Z(_11482_));
 OAI21_X2 _17358_ (.A(_10402_),
    .B1(_10344_),
    .B2(_10348_),
    .ZN(_11483_));
 AND2_X1 _17359_ (.A1(_10479_),
    .A2(_11483_),
    .ZN(_11484_));
 NAND3_X1 _17360_ (.A1(_11476_),
    .A2(_11482_),
    .A3(_11484_),
    .ZN(_11485_));
 BUF_X4 _17361_ (.A(_15362_),
    .Z(_11486_));
 NAND2_X4 _17362_ (.A1(_10479_),
    .A2(_11483_),
    .ZN(_11487_));
 OR3_X1 _17363_ (.A1(_11486_),
    .A2(_11481_),
    .A3(_11487_),
    .ZN(_11488_));
 OAI33_X1 _17364_ (.A1(_10340_),
    .A2(_10378_),
    .A3(_10554_),
    .B1(_11483_),
    .B2(_10368_),
    .B3(_10332_),
    .ZN(_11489_));
 OR2_X1 _17365_ (.A1(_10344_),
    .A2(_10482_),
    .ZN(_11490_));
 OAI21_X1 _17366_ (.A(_10483_),
    .B1(_10504_),
    .B2(_11490_),
    .ZN(_11491_));
 AOI211_X2 _17367_ (.A(_10533_),
    .B(net21),
    .C1(_11491_),
    .C2(_10487_),
    .ZN(_11492_));
 MUX2_X1 _17368_ (.A(net315),
    .B(_10347_),
    .S(_10670_),
    .Z(_11493_));
 NAND2_X1 _17369_ (.A1(_10508_),
    .A2(net282),
    .ZN(_11494_));
 OAI33_X1 _17370_ (.A1(_10347_),
    .A2(_10480_),
    .A3(_10481_),
    .B1(_10912_),
    .B2(_11494_),
    .B3(_10883_),
    .ZN(_11495_));
 NOR2_X2 _17371_ (.A1(_10380_),
    .A2(_10482_),
    .ZN(_11496_));
 AOI22_X4 _17372_ (.A1(_10479_),
    .A2(_11493_),
    .B1(_11496_),
    .B2(_11495_),
    .ZN(_11497_));
 OR3_X2 _17373_ (.A1(net315),
    .A2(_10490_),
    .A3(_10551_),
    .ZN(_11498_));
 AND2_X1 _17374_ (.A1(_10548_),
    .A2(_11498_),
    .ZN(_11499_));
 OAI211_X4 _17375_ (.A(_11492_),
    .B(_11497_),
    .C1(_10912_),
    .C2(_11499_),
    .ZN(_11500_));
 MUX2_X2 _17376_ (.A(_11485_),
    .B(_11488_),
    .S(_11500_),
    .Z(_11501_));
 NAND2_X1 _17377_ (.A1(_11405_),
    .A2(_11487_),
    .ZN(_11502_));
 INV_X1 _17378_ (.A(_15360_),
    .ZN(_11503_));
 AND2_X1 _17379_ (.A1(_11503_),
    .A2(_11481_),
    .ZN(_11504_));
 BUF_X4 _17380_ (.A(_15367_),
    .Z(_11505_));
 AND3_X1 _17381_ (.A1(_10333_),
    .A2(_10895_),
    .A3(_11493_),
    .ZN(_11506_));
 OAI33_X1 _17382_ (.A1(_10347_),
    .A2(_10480_),
    .A3(_10481_),
    .B1(_10512_),
    .B2(_10912_),
    .B3(_10498_),
    .ZN(_11507_));
 AOI21_X4 _17383_ (.A(_11506_),
    .B1(_11507_),
    .B2(_11496_),
    .ZN(_11508_));
 AND3_X1 _17384_ (.A1(_11505_),
    .A2(_11481_),
    .A3(_11508_),
    .ZN(_11509_));
 AOI21_X4 _17385_ (.A(_10912_),
    .B1(net277),
    .B2(_11498_),
    .ZN(_11510_));
 AND2_X1 _17386_ (.A1(_10487_),
    .A2(_11491_),
    .ZN(_11511_));
 NOR4_X4 _17387_ (.A1(_10533_),
    .A2(_11510_),
    .A3(_11511_),
    .A4(net21),
    .ZN(_11512_));
 MUX2_X2 _17388_ (.A(_11504_),
    .B(_11509_),
    .S(_11512_),
    .Z(_11513_));
 OAI21_X4 _17389_ (.A(_11501_),
    .B1(_11502_),
    .B2(_11513_),
    .ZN(_11514_));
 INV_X2 _17390_ (.A(_11514_),
    .ZN(_14064_));
 NOR3_X1 _17391_ (.A1(_00181_),
    .A2(_10565_),
    .A3(_10744_),
    .ZN(_11515_));
 AOI22_X2 _17392_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_10397_),
    .B1(_10683_),
    .B2(_11515_),
    .ZN(_11516_));
 BUF_X2 _17393_ (.A(\cs_registers_i.pc_id_i[3] ),
    .Z(_11517_));
 OAI21_X2 _17394_ (.A(_10565_),
    .B1(_10747_),
    .B2(_11517_),
    .ZN(_11518_));
 MUX2_X1 _17395_ (.A(_00285_),
    .B(_00287_),
    .S(_10588_),
    .Z(_11519_));
 MUX2_X1 _17396_ (.A(_00286_),
    .B(_00288_),
    .S(_10588_),
    .Z(_11520_));
 MUX2_X1 _17397_ (.A(_11519_),
    .B(_11520_),
    .S(_10629_),
    .Z(_11521_));
 NAND2_X1 _17398_ (.A1(_10767_),
    .A2(_11521_),
    .ZN(_11522_));
 NAND2_X1 _17399_ (.A1(_10616_),
    .A2(_00280_),
    .ZN(_11523_));
 OAI21_X1 _17400_ (.A(_11523_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .B2(_10616_),
    .ZN(_11524_));
 OAI221_X1 _17401_ (.A(_10571_),
    .B1(_00279_),
    .B2(_10758_),
    .C1(_11524_),
    .C2(_10582_),
    .ZN(_11525_));
 NAND4_X1 _17402_ (.A1(_10610_),
    .A2(_10576_),
    .A3(_11522_),
    .A4(_11525_),
    .ZN(_11526_));
 MUX2_X1 _17403_ (.A(_00297_),
    .B(_00299_),
    .S(_10600_),
    .Z(_11527_));
 MUX2_X1 _17404_ (.A(_00298_),
    .B(_00300_),
    .S(_10600_),
    .Z(_11528_));
 MUX2_X1 _17405_ (.A(_11527_),
    .B(_11528_),
    .S(_10628_),
    .Z(_11529_));
 MUX2_X1 _17406_ (.A(_00295_),
    .B(_00296_),
    .S(_10595_),
    .Z(_11530_));
 MUX2_X1 _17407_ (.A(_00293_),
    .B(_00294_),
    .S(_11366_),
    .Z(_11531_));
 AOI222_X2 _17408_ (.A1(_10778_),
    .A2(_11529_),
    .B1(_11530_),
    .B2(_10794_),
    .C1(_11531_),
    .C2(_10785_),
    .ZN(_11532_));
 BUF_X4 _17409_ (.A(_10766_),
    .Z(_11533_));
 BUF_X8 _17410_ (.A(_11383_),
    .Z(_11534_));
 BUF_X8 _17411_ (.A(_11534_),
    .Z(_11535_));
 MUX2_X1 _17412_ (.A(_00307_),
    .B(_00308_),
    .S(_11535_),
    .Z(_11536_));
 MUX2_X1 _17413_ (.A(_00305_),
    .B(_00306_),
    .S(_10797_),
    .Z(_11537_));
 OAI221_X1 _17414_ (.A(_11533_),
    .B1(_10838_),
    .B2(_11536_),
    .C1(_11537_),
    .C2(_10842_),
    .ZN(_11538_));
 MUX2_X1 _17415_ (.A(_00303_),
    .B(_00304_),
    .S(_10627_),
    .Z(_11539_));
 MUX2_X1 _17416_ (.A(_00301_),
    .B(_00302_),
    .S(_10787_),
    .Z(_11540_));
 MUX2_X1 _17417_ (.A(_11539_),
    .B(_11540_),
    .S(_10632_),
    .Z(_11541_));
 NOR2_X1 _17418_ (.A1(_10752_),
    .A2(_11541_),
    .ZN(_11542_));
 OAI21_X1 _17419_ (.A(_11532_),
    .B1(_11538_),
    .B2(_11542_),
    .ZN(_11543_));
 MUX2_X1 _17420_ (.A(_00289_),
    .B(_00291_),
    .S(_10614_),
    .Z(_11544_));
 BUF_X4 _17421_ (.A(_10857_),
    .Z(_11545_));
 BUF_X4 _17422_ (.A(_11545_),
    .Z(_11546_));
 BUF_X4 _17423_ (.A(_11546_),
    .Z(_11547_));
 MUX2_X1 _17424_ (.A(_00290_),
    .B(_00292_),
    .S(_11547_),
    .Z(_11548_));
 MUX2_X1 _17425_ (.A(_11544_),
    .B(_11548_),
    .S(_10596_),
    .Z(_11549_));
 MUX2_X1 _17426_ (.A(_00281_),
    .B(_00283_),
    .S(_11547_),
    .Z(_11550_));
 MUX2_X1 _17427_ (.A(_00282_),
    .B(_00284_),
    .S(_11547_),
    .Z(_11551_));
 MUX2_X1 _17428_ (.A(_11550_),
    .B(_11551_),
    .S(_10596_),
    .Z(_11552_));
 MUX2_X1 _17429_ (.A(_11549_),
    .B(_11552_),
    .S(_10570_),
    .Z(_11553_));
 OAI221_X2 _17430_ (.A(_11526_),
    .B1(_10576_),
    .B2(_11543_),
    .C1(_11553_),
    .C2(_10855_),
    .ZN(_11554_));
 NOR2_X1 _17431_ (.A1(_10683_),
    .A2(net319),
    .ZN(_11555_));
 OAI21_X4 _17432_ (.A(_11516_),
    .B1(_11518_),
    .B2(_11555_),
    .ZN(_15865_));
 INV_X2 _17433_ (.A(_15865_),
    .ZN(_15861_));
 INV_X1 _17434_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .ZN(_11556_));
 OR3_X2 _17435_ (.A1(_00180_),
    .A2(_10361_),
    .A3(_10743_),
    .ZN(_11557_));
 OAI22_X2 _17436_ (.A1(_11556_),
    .A2(_10673_),
    .B1(_10681_),
    .B2(_11557_),
    .ZN(_11558_));
 MUX2_X1 _17437_ (.A(_00323_),
    .B(_00325_),
    .S(_10600_),
    .Z(_11559_));
 MUX2_X1 _17438_ (.A(_00324_),
    .B(_00326_),
    .S(_10600_),
    .Z(_11560_));
 MUX2_X1 _17439_ (.A(_11559_),
    .B(_11560_),
    .S(_11535_),
    .Z(_11561_));
 AOI21_X1 _17440_ (.A(_11437_),
    .B1(_11561_),
    .B2(_11370_),
    .ZN(_11562_));
 NAND2_X1 _17441_ (.A1(_10621_),
    .A2(_00310_),
    .ZN(_11563_));
 OAI21_X1 _17442_ (.A(_11563_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B2(_10615_),
    .ZN(_11564_));
 OAI22_X1 _17443_ (.A1(_00309_),
    .A2(_10757_),
    .B1(_11564_),
    .B2(_10580_),
    .ZN(_11565_));
 OAI21_X2 _17444_ (.A(_11562_),
    .B1(_11565_),
    .B2(_10749_),
    .ZN(_11566_));
 BUF_X4 _17445_ (.A(_10611_),
    .Z(_11567_));
 BUF_X4 _17446_ (.A(_11567_),
    .Z(_11568_));
 MUX2_X1 _17447_ (.A(_00331_),
    .B(_00333_),
    .S(_11568_),
    .Z(_11569_));
 MUX2_X1 _17448_ (.A(_00332_),
    .B(_00334_),
    .S(_11568_),
    .Z(_11570_));
 MUX2_X1 _17449_ (.A(_11569_),
    .B(_11570_),
    .S(_10796_),
    .Z(_11571_));
 MUX2_X1 _17450_ (.A(_00315_),
    .B(_00317_),
    .S(_11568_),
    .Z(_11572_));
 MUX2_X1 _17451_ (.A(_00316_),
    .B(_00318_),
    .S(_11568_),
    .Z(_11573_));
 MUX2_X1 _17452_ (.A(_11572_),
    .B(_11573_),
    .S(_10796_),
    .Z(_11574_));
 MUX2_X1 _17453_ (.A(_11571_),
    .B(_11574_),
    .S(_10574_),
    .Z(_11575_));
 MUX2_X1 _17454_ (.A(_00335_),
    .B(_00337_),
    .S(_10618_),
    .Z(_11576_));
 MUX2_X1 _17455_ (.A(_00336_),
    .B(_00338_),
    .S(_10618_),
    .Z(_11577_));
 MUX2_X1 _17456_ (.A(_11576_),
    .B(_11577_),
    .S(_10795_),
    .Z(_11578_));
 MUX2_X1 _17457_ (.A(_00319_),
    .B(_00321_),
    .S(_10618_),
    .Z(_11579_));
 MUX2_X1 _17458_ (.A(_00320_),
    .B(_00322_),
    .S(_10618_),
    .Z(_11580_));
 MUX2_X1 _17459_ (.A(_11579_),
    .B(_11580_),
    .S(_10795_),
    .Z(_11581_));
 MUX2_X1 _17460_ (.A(_11578_),
    .B(_11581_),
    .S(_10573_),
    .Z(_11582_));
 MUX2_X1 _17461_ (.A(_00327_),
    .B(_00329_),
    .S(_10618_),
    .Z(_11583_));
 MUX2_X1 _17462_ (.A(_00328_),
    .B(_00330_),
    .S(_11567_),
    .Z(_11584_));
 MUX2_X1 _17463_ (.A(_11583_),
    .B(_11584_),
    .S(_10795_),
    .Z(_11585_));
 MUX2_X1 _17464_ (.A(_00311_),
    .B(_00313_),
    .S(_11567_),
    .Z(_11586_));
 MUX2_X1 _17465_ (.A(_00312_),
    .B(_00314_),
    .S(_11567_),
    .Z(_11587_));
 MUX2_X1 _17466_ (.A(_11586_),
    .B(_11587_),
    .S(_10795_),
    .Z(_11588_));
 MUX2_X1 _17467_ (.A(_11585_),
    .B(_11588_),
    .S(_10574_),
    .Z(_11589_));
 MUX2_X1 _17468_ (.A(_11582_),
    .B(_11589_),
    .S(_11358_),
    .Z(_11590_));
 OAI221_X2 _17469_ (.A(_11566_),
    .B1(_11575_),
    .B2(_11453_),
    .C1(_11590_),
    .C2(_10609_),
    .ZN(_11591_));
 AND2_X1 _17470_ (.A1(_10816_),
    .A2(_11591_),
    .ZN(_11592_));
 CLKBUF_X2 _17471_ (.A(_10563_),
    .Z(_11593_));
 AND2_X1 _17472_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_11593_),
    .ZN(_11594_));
 AND2_X1 _17473_ (.A1(_10683_),
    .A2(_11594_),
    .ZN(_11595_));
 OR3_X4 _17474_ (.A1(_11558_),
    .A2(_11592_),
    .A3(_11595_),
    .ZN(_15868_));
 INV_X2 _17475_ (.A(_15868_),
    .ZN(_15872_));
 BUF_X4 _17476_ (.A(_10816_),
    .Z(_11596_));
 BUF_X4 _17477_ (.A(_11568_),
    .Z(_11597_));
 MUX2_X1 _17478_ (.A(_00345_),
    .B(_00347_),
    .S(_11597_),
    .Z(_11598_));
 MUX2_X1 _17479_ (.A(_00346_),
    .B(_00348_),
    .S(_11597_),
    .Z(_11599_));
 MUX2_X1 _17480_ (.A(_11598_),
    .B(_11599_),
    .S(_10797_),
    .Z(_11600_));
 AOI21_X1 _17481_ (.A(_10831_),
    .B1(_11600_),
    .B2(_11533_),
    .ZN(_11601_));
 NAND2_X1 _17482_ (.A1(_10602_),
    .A2(_00340_),
    .ZN(_11602_));
 OAI21_X1 _17483_ (.A(_11602_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .B2(_10622_),
    .ZN(_11603_));
 OAI22_X1 _17484_ (.A1(_00339_),
    .A2(_10758_),
    .B1(_11603_),
    .B2(_10581_),
    .ZN(_11604_));
 OAI21_X1 _17485_ (.A(_11601_),
    .B1(_11604_),
    .B2(_10767_),
    .ZN(_11605_));
 MUX2_X1 _17486_ (.A(_00361_),
    .B(_00363_),
    .S(_11546_),
    .Z(_11606_));
 MUX2_X1 _17487_ (.A(_00362_),
    .B(_00364_),
    .S(_10823_),
    .Z(_11607_));
 MUX2_X1 _17488_ (.A(_11606_),
    .B(_11607_),
    .S(_11535_),
    .Z(_11608_));
 MUX2_X1 _17489_ (.A(_00353_),
    .B(_00355_),
    .S(_10823_),
    .Z(_11609_));
 MUX2_X1 _17490_ (.A(_00354_),
    .B(_00356_),
    .S(_10823_),
    .Z(_11610_));
 MUX2_X1 _17491_ (.A(_11609_),
    .B(_11610_),
    .S(_11535_),
    .Z(_11611_));
 MUX2_X1 _17492_ (.A(_11608_),
    .B(_11611_),
    .S(_11358_),
    .Z(_11612_));
 MUX2_X1 _17493_ (.A(_00365_),
    .B(_00367_),
    .S(_11545_),
    .Z(_11613_));
 BUF_X4 _17494_ (.A(_10598_),
    .Z(_11614_));
 MUX2_X1 _17495_ (.A(_00366_),
    .B(_00368_),
    .S(_11614_),
    .Z(_11615_));
 MUX2_X1 _17496_ (.A(_11613_),
    .B(_11615_),
    .S(_10594_),
    .Z(_11616_));
 MUX2_X1 _17497_ (.A(_00357_),
    .B(_00359_),
    .S(_11614_),
    .Z(_11617_));
 MUX2_X1 _17498_ (.A(_00358_),
    .B(_00360_),
    .S(_11614_),
    .Z(_11618_));
 MUX2_X1 _17499_ (.A(_11617_),
    .B(_11618_),
    .S(_10594_),
    .Z(_11619_));
 MUX2_X1 _17500_ (.A(_11616_),
    .B(_11619_),
    .S(_10569_),
    .Z(_11620_));
 MUX2_X1 _17501_ (.A(_00349_),
    .B(_00351_),
    .S(_11614_),
    .Z(_11621_));
 MUX2_X1 _17502_ (.A(_00350_),
    .B(_00352_),
    .S(_11614_),
    .Z(_11622_));
 MUX2_X1 _17503_ (.A(_11621_),
    .B(_11622_),
    .S(_10594_),
    .Z(_11623_));
 MUX2_X1 _17504_ (.A(_00341_),
    .B(_00343_),
    .S(_11614_),
    .Z(_11624_));
 MUX2_X1 _17505_ (.A(_00342_),
    .B(_00344_),
    .S(_11372_),
    .Z(_11625_));
 MUX2_X1 _17506_ (.A(_11624_),
    .B(_11625_),
    .S(_11375_),
    .Z(_11626_));
 MUX2_X1 _17507_ (.A(_11623_),
    .B(_11626_),
    .S(_10569_),
    .Z(_11627_));
 MUX2_X1 _17508_ (.A(_11620_),
    .B(_11627_),
    .S(_10783_),
    .Z(_11628_));
 OAI221_X2 _17509_ (.A(_11605_),
    .B1(_11612_),
    .B2(_11371_),
    .C1(_10609_),
    .C2(_11628_),
    .ZN(_11629_));
 AND2_X1 _17510_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_10564_),
    .ZN(_11630_));
 AOI222_X2 _17511_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(_10397_),
    .B1(_11596_),
    .B2(_11629_),
    .C1(_11630_),
    .C2(_10683_),
    .ZN(_11631_));
 BUF_X4 _17512_ (.A(_11631_),
    .Z(_15881_));
 BUF_X4 _17513_ (.A(_10361_),
    .Z(_11632_));
 MUX2_X1 _17514_ (.A(_00375_),
    .B(_00377_),
    .S(_10618_),
    .Z(_11633_));
 NOR2_X1 _17515_ (.A1(_10839_),
    .A2(_11633_),
    .ZN(_11634_));
 MUX2_X1 _17516_ (.A(_00376_),
    .B(_00378_),
    .S(_10618_),
    .Z(_11635_));
 NOR2_X1 _17517_ (.A1(_10579_),
    .A2(_11635_),
    .ZN(_11636_));
 NOR3_X1 _17518_ (.A1(_10568_),
    .A2(_11634_),
    .A3(_11636_),
    .ZN(_11637_));
 INV_X1 _17519_ (.A(_00369_),
    .ZN(_11638_));
 BUF_X4 _17520_ (.A(_10584_),
    .Z(_11639_));
 NOR2_X1 _17521_ (.A1(_11639_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .ZN(_11640_));
 BUF_X4 _17522_ (.A(_10856_),
    .Z(_11641_));
 BUF_X4 _17523_ (.A(_11641_),
    .Z(_11642_));
 AOI21_X1 _17524_ (.A(_11640_),
    .B1(_00370_),
    .B2(_11642_),
    .ZN(_11643_));
 AOI221_X2 _17525_ (.A(_10764_),
    .B1(_11638_),
    .B2(_10821_),
    .C1(_11643_),
    .C2(_11383_),
    .ZN(_11644_));
 NOR3_X2 _17526_ (.A1(_10832_),
    .A2(_11637_),
    .A3(_11644_),
    .ZN(_11645_));
 MUX2_X1 _17527_ (.A(_00379_),
    .B(_00381_),
    .S(_10611_),
    .Z(_11646_));
 MUX2_X1 _17528_ (.A(_00380_),
    .B(_00382_),
    .S(_10611_),
    .Z(_11647_));
 MUX2_X1 _17529_ (.A(_11646_),
    .B(_11647_),
    .S(_10625_),
    .Z(_11648_));
 MUX2_X1 _17530_ (.A(_00371_),
    .B(_00373_),
    .S(_10611_),
    .Z(_11649_));
 MUX2_X1 _17531_ (.A(_00372_),
    .B(_00374_),
    .S(_10611_),
    .Z(_11650_));
 MUX2_X1 _17532_ (.A(_11649_),
    .B(_11650_),
    .S(_10625_),
    .Z(_11651_));
 MUX2_X1 _17533_ (.A(_11648_),
    .B(_11651_),
    .S(_10567_),
    .Z(_11652_));
 NOR2_X1 _17534_ (.A1(_10607_),
    .A2(_11652_),
    .ZN(_11653_));
 NOR3_X2 _17535_ (.A1(_10572_),
    .A2(_11645_),
    .A3(_11653_),
    .ZN(_11654_));
 BUF_X4 _17536_ (.A(_10583_),
    .Z(_11655_));
 MUX2_X1 _17537_ (.A(_00391_),
    .B(_00393_),
    .S(_11655_),
    .Z(_11656_));
 MUX2_X1 _17538_ (.A(_00392_),
    .B(_00394_),
    .S(_11655_),
    .Z(_11657_));
 MUX2_X1 _17539_ (.A(_11656_),
    .B(_11657_),
    .S(_10833_),
    .Z(_11658_));
 MUX2_X1 _17540_ (.A(_00383_),
    .B(_00385_),
    .S(_11655_),
    .Z(_11659_));
 MUX2_X1 _17541_ (.A(_00384_),
    .B(_00386_),
    .S(_11655_),
    .Z(_11660_));
 MUX2_X1 _17542_ (.A(_11659_),
    .B(_11660_),
    .S(_10833_),
    .Z(_11661_));
 BUF_X4 _17543_ (.A(_10567_),
    .Z(_11662_));
 MUX2_X1 _17544_ (.A(_11658_),
    .B(_11661_),
    .S(_11662_),
    .Z(_11663_));
 MUX2_X1 _17545_ (.A(_00395_),
    .B(_00397_),
    .S(_11655_),
    .Z(_11664_));
 MUX2_X1 _17546_ (.A(_00396_),
    .B(_00398_),
    .S(_10790_),
    .Z(_11665_));
 MUX2_X1 _17547_ (.A(_11664_),
    .B(_11665_),
    .S(_10833_),
    .Z(_11666_));
 MUX2_X1 _17548_ (.A(_00387_),
    .B(_00389_),
    .S(_10790_),
    .Z(_11667_));
 MUX2_X1 _17549_ (.A(_00388_),
    .B(_00390_),
    .S(_10790_),
    .Z(_11668_));
 MUX2_X1 _17550_ (.A(_11667_),
    .B(_11668_),
    .S(_10833_),
    .Z(_11669_));
 MUX2_X1 _17551_ (.A(_11666_),
    .B(_11669_),
    .S(_11662_),
    .Z(_11670_));
 MUX2_X1 _17552_ (.A(_11663_),
    .B(_11670_),
    .S(_10832_),
    .Z(_11671_));
 AOI21_X4 _17553_ (.A(_11654_),
    .B1(_11671_),
    .B2(_11370_),
    .ZN(_11672_));
 INV_X1 _17554_ (.A(\cs_registers_i.pc_id_i[6] ),
    .ZN(_11673_));
 NOR2_X1 _17555_ (.A1(_11673_),
    .A2(_10668_),
    .ZN(_11674_));
 AOI222_X2 _17556_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(_11632_),
    .B1(_10816_),
    .B2(_11672_),
    .C1(_11674_),
    .C2(_10682_),
    .ZN(_15889_));
 NAND2_X1 _17557_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(_11632_),
    .ZN(_11675_));
 BUF_X4 _17558_ (.A(_10606_),
    .Z(_11676_));
 MUX2_X1 _17559_ (.A(_00421_),
    .B(_00423_),
    .S(_11639_),
    .Z(_11677_));
 BUF_X4 _17560_ (.A(_10584_),
    .Z(_11678_));
 MUX2_X1 _17561_ (.A(_00422_),
    .B(_00424_),
    .S(_11678_),
    .Z(_11679_));
 MUX2_X1 _17562_ (.A(_11677_),
    .B(_11679_),
    .S(_10626_),
    .Z(_11680_));
 MUX2_X1 _17563_ (.A(_00413_),
    .B(_00415_),
    .S(_11678_),
    .Z(_11681_));
 MUX2_X1 _17564_ (.A(_00414_),
    .B(_00416_),
    .S(_11678_),
    .Z(_11682_));
 MUX2_X1 _17565_ (.A(_11681_),
    .B(_11682_),
    .S(_10626_),
    .Z(_11683_));
 MUX2_X1 _17566_ (.A(_11680_),
    .B(_11683_),
    .S(_10827_),
    .Z(_11684_));
 NOR2_X2 _17567_ (.A1(_11676_),
    .A2(_11684_),
    .ZN(_11685_));
 MUX2_X1 _17568_ (.A(_00425_),
    .B(_00427_),
    .S(_11639_),
    .Z(_11686_));
 MUX2_X1 _17569_ (.A(_00426_),
    .B(_00428_),
    .S(_11639_),
    .Z(_11687_));
 MUX2_X1 _17570_ (.A(_11686_),
    .B(_11687_),
    .S(_10626_),
    .Z(_11688_));
 MUX2_X1 _17571_ (.A(_00417_),
    .B(_00419_),
    .S(_11639_),
    .Z(_11689_));
 MUX2_X1 _17572_ (.A(_00418_),
    .B(_00420_),
    .S(_11639_),
    .Z(_11690_));
 MUX2_X1 _17573_ (.A(_11689_),
    .B(_11690_),
    .S(_10626_),
    .Z(_11691_));
 MUX2_X1 _17574_ (.A(_11688_),
    .B(_11691_),
    .S(_10568_),
    .Z(_11692_));
 NOR2_X1 _17575_ (.A1(_10608_),
    .A2(_11692_),
    .ZN(_11693_));
 NOR3_X4 _17576_ (.A1(_10783_),
    .A2(_11685_),
    .A3(_11693_),
    .ZN(_11694_));
 MUX2_X1 _17577_ (.A(_00405_),
    .B(_00407_),
    .S(_10599_),
    .Z(_11695_));
 NOR2_X1 _17578_ (.A1(_10796_),
    .A2(_11695_),
    .ZN(_11696_));
 MUX2_X1 _17579_ (.A(_00406_),
    .B(_00408_),
    .S(_11372_),
    .Z(_11697_));
 NOR2_X1 _17580_ (.A1(_10579_),
    .A2(_11697_),
    .ZN(_11698_));
 NOR3_X1 _17581_ (.A1(_11357_),
    .A2(_11696_),
    .A3(_11698_),
    .ZN(_11699_));
 INV_X1 _17582_ (.A(_00399_),
    .ZN(_11700_));
 NOR2_X1 _17583_ (.A1(_11642_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .ZN(_11701_));
 AOI21_X1 _17584_ (.A(_11701_),
    .B1(_00400_),
    .B2(_11568_),
    .ZN(_11702_));
 AOI221_X2 _17585_ (.A(_10765_),
    .B1(_11700_),
    .B2(_10822_),
    .C1(_11702_),
    .C2(_10839_),
    .ZN(_11703_));
 NOR3_X2 _17586_ (.A1(_11676_),
    .A2(_11699_),
    .A3(_11703_),
    .ZN(_11704_));
 MUX2_X1 _17587_ (.A(_00409_),
    .B(_00411_),
    .S(_10598_),
    .Z(_11705_));
 MUX2_X1 _17588_ (.A(_00410_),
    .B(_00412_),
    .S(_10598_),
    .Z(_11706_));
 MUX2_X1 _17589_ (.A(_11705_),
    .B(_11706_),
    .S(_11383_),
    .Z(_11707_));
 MUX2_X1 _17590_ (.A(_00401_),
    .B(_00403_),
    .S(_10598_),
    .Z(_11708_));
 MUX2_X1 _17591_ (.A(_00402_),
    .B(_00404_),
    .S(_10598_),
    .Z(_11709_));
 MUX2_X1 _17592_ (.A(_11708_),
    .B(_11709_),
    .S(_11383_),
    .Z(_11710_));
 MUX2_X1 _17593_ (.A(_11707_),
    .B(_11710_),
    .S(_10568_),
    .Z(_11711_));
 NOR2_X2 _17594_ (.A1(_10608_),
    .A2(_11711_),
    .ZN(_11712_));
 NOR3_X4 _17595_ (.A1(_11370_),
    .A2(_11704_),
    .A3(_11712_),
    .ZN(_11713_));
 OR2_X2 _17596_ (.A1(_11694_),
    .A2(_11713_),
    .ZN(_11714_));
 NAND2_X1 _17597_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_10564_),
    .ZN(_11715_));
 OAI221_X1 _17598_ (.A(_11675_),
    .B1(_11714_),
    .B2(_10814_),
    .C1(_11715_),
    .C2(_10747_),
    .ZN(_11716_));
 CLKBUF_X3 _17599_ (.A(_11716_),
    .Z(_15893_));
 INV_X1 _17600_ (.A(_15893_),
    .ZN(_15897_));
 BUF_X2 _17601_ (.A(_15398_),
    .Z(_11717_));
 INV_X1 _17602_ (.A(_15385_),
    .ZN(_11718_));
 AOI21_X2 _17603_ (.A(_15371_),
    .B1(_14067_),
    .B2(_10815_),
    .ZN(_11719_));
 BUF_X2 _17604_ (.A(_15378_),
    .Z(_11720_));
 BUF_X4 _17605_ (.A(_15382_),
    .Z(_11721_));
 BUF_X2 _17606_ (.A(_15386_),
    .Z(_11722_));
 NAND3_X1 _17607_ (.A1(_11720_),
    .A2(_11721_),
    .A3(_11722_),
    .ZN(_11723_));
 AOI21_X2 _17608_ (.A(_15381_),
    .B1(_15377_),
    .B2(_11721_),
    .ZN(_11724_));
 INV_X1 _17609_ (.A(_11722_),
    .ZN(_11725_));
 OAI221_X2 _17610_ (.A(_11718_),
    .B1(_11723_),
    .B2(_11719_),
    .C1(_11724_),
    .C2(_11725_),
    .ZN(_11726_));
 BUF_X1 _17611_ (.A(_15390_),
    .Z(_11727_));
 AOI21_X1 _17612_ (.A(_15389_),
    .B1(_11726_),
    .B2(_11727_),
    .ZN(_11728_));
 INV_X1 _17613_ (.A(_11728_),
    .ZN(_11729_));
 BUF_X2 _17614_ (.A(_15394_),
    .Z(_11730_));
 AOI21_X2 _17615_ (.A(_15393_),
    .B1(_11729_),
    .B2(_11730_),
    .ZN(_11731_));
 XNOR2_X2 _17616_ (.A(_11717_),
    .B(_11731_),
    .ZN(\alu_adder_result_ex[7] ));
 INV_X1 _17617_ (.A(_15389_),
    .ZN(_11732_));
 INV_X1 _17618_ (.A(_11724_),
    .ZN(_11733_));
 AOI21_X1 _17619_ (.A(_15385_),
    .B1(_11733_),
    .B2(_11722_),
    .ZN(_11734_));
 INV_X1 _17620_ (.A(_11727_),
    .ZN(_11735_));
 OAI21_X1 _17621_ (.A(_11732_),
    .B1(_11734_),
    .B2(_11735_),
    .ZN(_11736_));
 NAND2_X2 _17622_ (.A1(_11720_),
    .A2(_11721_),
    .ZN(_11737_));
 NAND2_X1 _17623_ (.A1(_11722_),
    .A2(_11727_),
    .ZN(_11738_));
 AOI21_X2 _17624_ (.A(_15371_),
    .B1(_15373_),
    .B2(_10815_),
    .ZN(_11739_));
 NOR3_X1 _17625_ (.A1(_11737_),
    .A2(_11738_),
    .A3(_11739_),
    .ZN(_11740_));
 NOR2_X1 _17626_ (.A1(_11736_),
    .A2(_11740_),
    .ZN(_11741_));
 XNOR2_X1 _17627_ (.A(_11730_),
    .B(_11741_),
    .ZN(_11742_));
 NOR2_X1 _17628_ (.A1(_11737_),
    .A2(_11738_),
    .ZN(_11743_));
 NAND2_X4 _17629_ (.A1(_15374_),
    .A2(_10815_),
    .ZN(_11744_));
 NAND2_X1 _17630_ (.A1(_11739_),
    .A2(_11744_),
    .ZN(_11745_));
 AOI21_X1 _17631_ (.A(_11736_),
    .B1(_11743_),
    .B2(_11745_),
    .ZN(_11746_));
 XNOR2_X1 _17632_ (.A(_11730_),
    .B(_11746_),
    .ZN(_11747_));
 MUX2_X1 _17633_ (.A(_11742_),
    .B(_11747_),
    .S(_14064_),
    .Z(_11748_));
 BUF_X4 _17634_ (.A(_11748_),
    .Z(\alu_adder_result_ex[6] ));
 NAND2_X1 _17635_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(_11632_),
    .ZN(_11749_));
 MUX2_X1 _17636_ (.A(_00455_),
    .B(_00457_),
    .S(_10585_),
    .Z(_11750_));
 MUX2_X1 _17637_ (.A(_00456_),
    .B(_00458_),
    .S(_10585_),
    .Z(_11751_));
 MUX2_X1 _17638_ (.A(_11750_),
    .B(_11751_),
    .S(_10786_),
    .Z(_11752_));
 MUX2_X1 _17639_ (.A(_00447_),
    .B(_00449_),
    .S(_10585_),
    .Z(_11753_));
 MUX2_X1 _17640_ (.A(_00448_),
    .B(_00450_),
    .S(_10585_),
    .Z(_11754_));
 MUX2_X1 _17641_ (.A(_11753_),
    .B(_11754_),
    .S(_10786_),
    .Z(_11755_));
 MUX2_X1 _17642_ (.A(_11752_),
    .B(_11755_),
    .S(_10827_),
    .Z(_11756_));
 NAND2_X1 _17643_ (.A1(_11676_),
    .A2(_11756_),
    .ZN(_11757_));
 MUX2_X1 _17644_ (.A(_00451_),
    .B(_00453_),
    .S(_11545_),
    .Z(_11758_));
 MUX2_X1 _17645_ (.A(_00452_),
    .B(_00454_),
    .S(_11545_),
    .Z(_11759_));
 MUX2_X1 _17646_ (.A(_11758_),
    .B(_11759_),
    .S(_10594_),
    .Z(_11760_));
 MUX2_X1 _17647_ (.A(_00445_),
    .B(_00446_),
    .S(_10843_),
    .Z(_11761_));
 MUX2_X1 _17648_ (.A(_00443_),
    .B(_00444_),
    .S(_10795_),
    .Z(_11762_));
 AOI222_X2 _17649_ (.A1(_10643_),
    .A2(_11760_),
    .B1(_11761_),
    .B2(_10794_),
    .C1(_11762_),
    .C2(_10785_),
    .ZN(_11763_));
 AOI21_X4 _17650_ (.A(_10783_),
    .B1(_11757_),
    .B2(_11763_),
    .ZN(_11764_));
 MUX2_X1 _17651_ (.A(_00435_),
    .B(_00437_),
    .S(_11362_),
    .Z(_11765_));
 NOR2_X1 _17652_ (.A1(_11534_),
    .A2(_11765_),
    .ZN(_11766_));
 MUX2_X1 _17653_ (.A(_00436_),
    .B(_00438_),
    .S(_11362_),
    .Z(_11767_));
 NOR2_X1 _17654_ (.A1(_10579_),
    .A2(_11767_),
    .ZN(_11768_));
 NOR3_X1 _17655_ (.A1(_10827_),
    .A2(_11766_),
    .A3(_11768_),
    .ZN(_11769_));
 NOR2_X1 _17656_ (.A1(_11567_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .ZN(_11770_));
 BUF_X4 _17657_ (.A(_11639_),
    .Z(_11771_));
 AOI21_X1 _17658_ (.A(_11770_),
    .B1(_00430_),
    .B2(_11771_),
    .ZN(_11772_));
 AOI221_X2 _17659_ (.A(_10765_),
    .B1(_11226_),
    .B2(_10822_),
    .C1(_11772_),
    .C2(_10795_),
    .ZN(_11773_));
 NOR3_X2 _17660_ (.A1(_10832_),
    .A2(_11769_),
    .A3(_11773_),
    .ZN(_11774_));
 BUF_X4 _17661_ (.A(_10607_),
    .Z(_11775_));
 BUF_X4 _17662_ (.A(_10856_),
    .Z(_11776_));
 MUX2_X1 _17663_ (.A(_00439_),
    .B(_00441_),
    .S(_11776_),
    .Z(_11777_));
 BUF_X4 _17664_ (.A(_10856_),
    .Z(_11778_));
 MUX2_X1 _17665_ (.A(_00440_),
    .B(_00442_),
    .S(_11778_),
    .Z(_11779_));
 MUX2_X1 _17666_ (.A(_11777_),
    .B(_11779_),
    .S(_10839_),
    .Z(_11780_));
 MUX2_X1 _17667_ (.A(_00431_),
    .B(_00433_),
    .S(_11778_),
    .Z(_11781_));
 MUX2_X1 _17668_ (.A(_00432_),
    .B(_00434_),
    .S(_11778_),
    .Z(_11782_));
 MUX2_X1 _17669_ (.A(_11781_),
    .B(_11782_),
    .S(_10839_),
    .Z(_11783_));
 MUX2_X1 _17670_ (.A(_11780_),
    .B(_11783_),
    .S(_11662_),
    .Z(_11784_));
 NOR2_X1 _17671_ (.A1(_11775_),
    .A2(_11784_),
    .ZN(_11785_));
 NOR3_X4 _17672_ (.A1(_11370_),
    .A2(_11774_),
    .A3(_11785_),
    .ZN(_11786_));
 OR2_X2 _17673_ (.A1(_11764_),
    .A2(_11786_),
    .ZN(_11787_));
 CLKBUF_X2 _17674_ (.A(\cs_registers_i.pc_id_i[8] ),
    .Z(_11788_));
 NAND2_X1 _17675_ (.A1(_11788_),
    .A2(_10564_),
    .ZN(_11789_));
 OAI221_X2 _17676_ (.A(_11749_),
    .B1(_11787_),
    .B2(_10814_),
    .C1(_11789_),
    .C2(_10747_),
    .ZN(_15901_));
 INV_X2 _17677_ (.A(_15901_),
    .ZN(_15905_));
 NAND2_X1 _17678_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(_11632_),
    .ZN(_11790_));
 MUX2_X1 _17679_ (.A(_00465_),
    .B(_00467_),
    .S(_11567_),
    .Z(_11791_));
 NOR2_X1 _17680_ (.A1(_10862_),
    .A2(_11791_),
    .ZN(_11792_));
 MUX2_X1 _17681_ (.A(_00466_),
    .B(_00468_),
    .S(_10618_),
    .Z(_11793_));
 NOR2_X1 _17682_ (.A1(_10579_),
    .A2(_11793_),
    .ZN(_11794_));
 NOR3_X1 _17683_ (.A1(_10568_),
    .A2(_11792_),
    .A3(_11794_),
    .ZN(_11795_));
 NOR2_X1 _17684_ (.A1(_11639_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .ZN(_11796_));
 AOI21_X1 _17685_ (.A(_11796_),
    .B1(_00460_),
    .B2(_11642_),
    .ZN(_11797_));
 AOI221_X1 _17686_ (.A(_10764_),
    .B1(_11273_),
    .B2(_10821_),
    .C1(_11797_),
    .C2(_10626_),
    .ZN(_11798_));
 NOR3_X1 _17687_ (.A1(_10832_),
    .A2(_11795_),
    .A3(_11798_),
    .ZN(_11799_));
 MUX2_X1 _17688_ (.A(_00469_),
    .B(_00471_),
    .S(_10611_),
    .Z(_11800_));
 MUX2_X1 _17689_ (.A(_00470_),
    .B(_00472_),
    .S(_10611_),
    .Z(_11801_));
 MUX2_X1 _17690_ (.A(_11800_),
    .B(_11801_),
    .S(_10625_),
    .Z(_11802_));
 MUX2_X1 _17691_ (.A(_00461_),
    .B(_00463_),
    .S(_10611_),
    .Z(_11803_));
 MUX2_X1 _17692_ (.A(_00462_),
    .B(_00464_),
    .S(_10611_),
    .Z(_11804_));
 MUX2_X1 _17693_ (.A(_11803_),
    .B(_11804_),
    .S(_10625_),
    .Z(_11805_));
 MUX2_X1 _17694_ (.A(_11802_),
    .B(_11805_),
    .S(_10567_),
    .Z(_11806_));
 NOR2_X1 _17695_ (.A1(_11775_),
    .A2(_11806_),
    .ZN(_11807_));
 NOR3_X2 _17696_ (.A1(_11370_),
    .A2(_11799_),
    .A3(_11807_),
    .ZN(_11808_));
 MUX2_X1 _17697_ (.A(_00481_),
    .B(_00483_),
    .S(_11776_),
    .Z(_11809_));
 MUX2_X1 _17698_ (.A(_00482_),
    .B(_00484_),
    .S(_11776_),
    .Z(_11810_));
 MUX2_X1 _17699_ (.A(_11809_),
    .B(_11810_),
    .S(_10839_),
    .Z(_11811_));
 MUX2_X1 _17700_ (.A(_00473_),
    .B(_00475_),
    .S(_11776_),
    .Z(_11812_));
 MUX2_X1 _17701_ (.A(_00474_),
    .B(_00476_),
    .S(_11776_),
    .Z(_11813_));
 MUX2_X1 _17702_ (.A(_11812_),
    .B(_11813_),
    .S(_10839_),
    .Z(_11814_));
 MUX2_X1 _17703_ (.A(_11811_),
    .B(_11814_),
    .S(_11662_),
    .Z(_11815_));
 MUX2_X1 _17704_ (.A(_00485_),
    .B(_00487_),
    .S(_11776_),
    .Z(_11816_));
 MUX2_X1 _17705_ (.A(_00486_),
    .B(_00488_),
    .S(_11778_),
    .Z(_11817_));
 MUX2_X1 _17706_ (.A(_11816_),
    .B(_11817_),
    .S(_10839_),
    .Z(_11818_));
 MUX2_X1 _17707_ (.A(_00477_),
    .B(_00479_),
    .S(_11776_),
    .Z(_11819_));
 MUX2_X1 _17708_ (.A(_00478_),
    .B(_00480_),
    .S(_11778_),
    .Z(_11820_));
 MUX2_X1 _17709_ (.A(_11819_),
    .B(_11820_),
    .S(_10839_),
    .Z(_11821_));
 MUX2_X1 _17710_ (.A(_11818_),
    .B(_11821_),
    .S(_11662_),
    .Z(_11822_));
 MUX2_X1 _17711_ (.A(_11815_),
    .B(_11822_),
    .S(_10832_),
    .Z(_11823_));
 AOI21_X4 _17712_ (.A(_11808_),
    .B1(_11823_),
    .B2(_10749_),
    .ZN(_11824_));
 INV_X1 _17713_ (.A(_11824_),
    .ZN(_11825_));
 BUF_X1 _17714_ (.A(\cs_registers_i.pc_id_i[9] ),
    .Z(_11826_));
 NAND2_X1 _17715_ (.A1(_11826_),
    .A2(_10564_),
    .ZN(_11827_));
 OAI221_X2 _17716_ (.A(_11790_),
    .B1(_11825_),
    .B2(_10814_),
    .C1(_11827_),
    .C2(_10747_),
    .ZN(_15909_));
 INV_X2 _17717_ (.A(_15909_),
    .ZN(_15913_));
 BUF_X2 _17718_ (.A(_15406_),
    .Z(_11828_));
 INV_X1 _17719_ (.A(_15401_),
    .ZN(_11829_));
 AND3_X1 _17720_ (.A1(_11717_),
    .A2(_11727_),
    .A3(_11730_),
    .ZN(_11830_));
 AOI21_X1 _17721_ (.A(_15393_),
    .B1(_15389_),
    .B2(_11730_),
    .ZN(_11831_));
 INV_X1 _17722_ (.A(_11831_),
    .ZN(_11832_));
 AOI221_X2 _17723_ (.A(_15397_),
    .B1(_11726_),
    .B2(_11830_),
    .C1(_11832_),
    .C2(_11717_),
    .ZN(_11833_));
 BUF_X2 _17724_ (.A(_15402_),
    .Z(_11834_));
 INV_X1 _17725_ (.A(_11834_),
    .ZN(_11835_));
 OAI21_X1 _17726_ (.A(_11829_),
    .B1(_11833_),
    .B2(_11835_),
    .ZN(_11836_));
 XOR2_X2 _17727_ (.A(_11836_),
    .B(_11828_),
    .Z(\alu_adder_result_ex[9] ));
 AND2_X1 _17728_ (.A1(_11717_),
    .A2(_11730_),
    .ZN(_11837_));
 NOR2_X4 _17729_ (.A1(_11737_),
    .A2(_11744_),
    .ZN(_11838_));
 AND4_X4 _17730_ (.A1(_11722_),
    .A2(_11727_),
    .A3(_11837_),
    .A4(_11838_),
    .ZN(_11839_));
 NOR2_X1 _17731_ (.A1(_11834_),
    .A2(_11839_),
    .ZN(_11840_));
 INV_X1 _17732_ (.A(_15377_),
    .ZN(_11841_));
 INV_X1 _17733_ (.A(_11720_),
    .ZN(_11842_));
 OAI21_X1 _17734_ (.A(_11841_),
    .B1(_11739_),
    .B2(_11842_),
    .ZN(_11843_));
 AOI21_X2 _17735_ (.A(_15381_),
    .B1(_11843_),
    .B2(_11721_),
    .ZN(_11844_));
 NAND4_X1 _17736_ (.A1(_10873_),
    .A2(_10514_),
    .A3(_10917_),
    .A4(_11838_),
    .ZN(_11845_));
 AOI21_X2 _17737_ (.A(_11738_),
    .B1(_11844_),
    .B2(_11845_),
    .ZN(_11846_));
 OAI21_X2 _17738_ (.A(_11732_),
    .B1(_11718_),
    .B2(_11735_),
    .ZN(_11847_));
 OAI21_X4 _17739_ (.A(_11837_),
    .B1(_11846_),
    .B2(_11847_),
    .ZN(_11848_));
 AOI21_X2 _17740_ (.A(_15397_),
    .B1(_15393_),
    .B2(_11717_),
    .ZN(_11849_));
 AND2_X1 _17741_ (.A1(_11848_),
    .A2(_11849_),
    .ZN(_11850_));
 MUX2_X1 _17742_ (.A(_11834_),
    .B(_11840_),
    .S(_11850_),
    .Z(_11851_));
 AND3_X1 _17743_ (.A1(_11476_),
    .A2(_11482_),
    .A3(_11484_),
    .ZN(_11852_));
 NOR3_X1 _17744_ (.A1(_11486_),
    .A2(_11482_),
    .A3(_11487_),
    .ZN(_11853_));
 MUX2_X2 _17745_ (.A(_11852_),
    .B(_11853_),
    .S(_11500_),
    .Z(_11854_));
 NAND2_X1 _17746_ (.A1(_11834_),
    .A2(_11839_),
    .ZN(_11855_));
 NAND2_X1 _17747_ (.A1(_11503_),
    .A2(_11482_),
    .ZN(_11856_));
 NAND3_X2 _17748_ (.A1(_11505_),
    .A2(_11482_),
    .A3(_11508_),
    .ZN(_11857_));
 MUX2_X2 _17749_ (.A(_11856_),
    .B(_11857_),
    .S(_11512_),
    .Z(_11858_));
 AOI211_X2 _17750_ (.A(_11854_),
    .B(_11855_),
    .C1(_11858_),
    .C2(_11487_),
    .ZN(_11859_));
 NAND2_X2 _17751_ (.A1(_11848_),
    .A2(_11849_),
    .ZN(_11860_));
 NOR2_X1 _17752_ (.A1(_11834_),
    .A2(_11860_),
    .ZN(_11861_));
 BUF_X4 _17753_ (.A(_11484_),
    .Z(_11862_));
 OAI21_X4 _17754_ (.A(_11501_),
    .B1(_11862_),
    .B2(_11513_),
    .ZN(_11863_));
 AOI211_X4 _17755_ (.A(_11851_),
    .B(_11859_),
    .C1(_11861_),
    .C2(_11863_),
    .ZN(\alu_adder_result_ex[8] ));
 AND2_X1 _17756_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(_11593_),
    .ZN(_11864_));
 AOI22_X2 _17757_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(_10741_),
    .B1(_10870_),
    .B2(_11864_),
    .ZN(_11865_));
 MUX2_X1 _17758_ (.A(_00495_),
    .B(_00497_),
    .S(_10587_),
    .Z(_11866_));
 MUX2_X1 _17759_ (.A(_00496_),
    .B(_00498_),
    .S(_10587_),
    .Z(_11867_));
 MUX2_X1 _17760_ (.A(_11866_),
    .B(_11867_),
    .S(_10788_),
    .Z(_11868_));
 AOI21_X1 _17761_ (.A(_10831_),
    .B1(_11868_),
    .B2(_10766_),
    .ZN(_11869_));
 NAND2_X1 _17762_ (.A1(_10615_),
    .A2(_00490_),
    .ZN(_11870_));
 OAI21_X1 _17763_ (.A(_11870_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .B2(_10589_),
    .ZN(_11871_));
 OAI22_X1 _17764_ (.A1(_00489_),
    .A2(_10758_),
    .B1(_11871_),
    .B2(_10581_),
    .ZN(_11872_));
 OAI21_X1 _17765_ (.A(_11869_),
    .B1(_11872_),
    .B2(_11533_),
    .ZN(_11873_));
 BUF_X4 _17766_ (.A(_11362_),
    .Z(_11874_));
 MUX2_X1 _17767_ (.A(_00511_),
    .B(_00513_),
    .S(_11874_),
    .Z(_11875_));
 MUX2_X1 _17768_ (.A(_00512_),
    .B(_00514_),
    .S(_11363_),
    .Z(_11876_));
 BUF_X4 _17769_ (.A(_10843_),
    .Z(_11877_));
 MUX2_X1 _17770_ (.A(_11875_),
    .B(_11876_),
    .S(_11877_),
    .Z(_11878_));
 MUX2_X1 _17771_ (.A(_00503_),
    .B(_00505_),
    .S(_11363_),
    .Z(_11879_));
 MUX2_X1 _17772_ (.A(_00504_),
    .B(_00506_),
    .S(_11363_),
    .Z(_11880_));
 MUX2_X1 _17773_ (.A(_11879_),
    .B(_11880_),
    .S(_11366_),
    .Z(_11881_));
 MUX2_X1 _17774_ (.A(_11878_),
    .B(_11881_),
    .S(_11358_),
    .Z(_11882_));
 MUX2_X1 _17775_ (.A(_00515_),
    .B(_00517_),
    .S(_10791_),
    .Z(_11883_));
 MUX2_X1 _17776_ (.A(_00516_),
    .B(_00518_),
    .S(_10791_),
    .Z(_11884_));
 MUX2_X1 _17777_ (.A(_11883_),
    .B(_11884_),
    .S(_10839_),
    .Z(_11885_));
 MUX2_X1 _17778_ (.A(_00507_),
    .B(_00509_),
    .S(_10791_),
    .Z(_11886_));
 MUX2_X1 _17779_ (.A(_00508_),
    .B(_00510_),
    .S(_10791_),
    .Z(_11887_));
 MUX2_X1 _17780_ (.A(_11886_),
    .B(_11887_),
    .S(_10839_),
    .Z(_11888_));
 MUX2_X1 _17781_ (.A(_11885_),
    .B(_11888_),
    .S(_11357_),
    .Z(_11889_));
 MUX2_X1 _17782_ (.A(_00499_),
    .B(_00501_),
    .S(_10791_),
    .Z(_11890_));
 MUX2_X1 _17783_ (.A(_00500_),
    .B(_00502_),
    .S(_10791_),
    .Z(_11891_));
 MUX2_X1 _17784_ (.A(_11890_),
    .B(_11891_),
    .S(_10839_),
    .Z(_11892_));
 MUX2_X1 _17785_ (.A(_00491_),
    .B(_00493_),
    .S(_10791_),
    .Z(_11893_));
 MUX2_X1 _17786_ (.A(_00492_),
    .B(_00494_),
    .S(_10791_),
    .Z(_11894_));
 MUX2_X1 _17787_ (.A(_11893_),
    .B(_11894_),
    .S(_10839_),
    .Z(_11895_));
 MUX2_X1 _17788_ (.A(_11892_),
    .B(_11895_),
    .S(_11357_),
    .Z(_11896_));
 MUX2_X1 _17789_ (.A(_11889_),
    .B(_11896_),
    .S(_10575_),
    .Z(_11897_));
 OAI221_X2 _17790_ (.A(_11873_),
    .B1(_11882_),
    .B2(_11371_),
    .C1(_10609_),
    .C2(_11897_),
    .ZN(_11898_));
 INV_X1 _17791_ (.A(_11898_),
    .ZN(_11899_));
 OAI21_X2 _17792_ (.A(_11865_),
    .B1(_11899_),
    .B2(_10814_),
    .ZN(_15917_));
 INV_X2 _17793_ (.A(_15917_),
    .ZN(_15921_));
 BUF_X2 _17794_ (.A(_15414_),
    .Z(_11900_));
 CLKBUF_X2 _17795_ (.A(_15409_),
    .Z(_11901_));
 CLKBUF_X2 _17796_ (.A(_15410_),
    .Z(_11902_));
 INV_X1 _17797_ (.A(_11902_),
    .ZN(_11903_));
 AOI21_X2 _17798_ (.A(_15405_),
    .B1(_15401_),
    .B2(_11828_),
    .ZN(_11904_));
 NAND2_X2 _17799_ (.A1(_11834_),
    .A2(_11828_),
    .ZN(_11905_));
 AOI21_X1 _17800_ (.A(_11903_),
    .B1(_11904_),
    .B2(_11905_),
    .ZN(_11906_));
 OAI21_X2 _17801_ (.A(_11900_),
    .B1(_11901_),
    .B2(_11906_),
    .ZN(_11907_));
 INV_X1 _17802_ (.A(_11901_),
    .ZN(_11908_));
 AND2_X1 _17803_ (.A1(_11908_),
    .A2(_11904_),
    .ZN(_11909_));
 AOI21_X4 _17804_ (.A(_11907_),
    .B1(_11833_),
    .B2(_11909_),
    .ZN(_11910_));
 NOR2_X1 _17805_ (.A1(_11900_),
    .A2(_11901_),
    .ZN(_11911_));
 OAI21_X1 _17806_ (.A(_11904_),
    .B1(_11905_),
    .B2(_11833_),
    .ZN(_11912_));
 NAND2_X1 _17807_ (.A1(_11902_),
    .A2(_11912_),
    .ZN(_11913_));
 AOI21_X4 _17808_ (.A(_11910_),
    .B1(_11911_),
    .B2(_11913_),
    .ZN(\alu_adder_result_ex[11] ));
 OAI21_X1 _17809_ (.A(_11829_),
    .B1(_11849_),
    .B2(_11835_),
    .ZN(_11914_));
 AOI21_X2 _17810_ (.A(_15405_),
    .B1(_11914_),
    .B2(_11828_),
    .ZN(_11915_));
 OAI21_X4 _17811_ (.A(_11915_),
    .B1(_11905_),
    .B2(_11848_),
    .ZN(_11916_));
 NAND3_X1 _17812_ (.A1(_11834_),
    .A2(_11828_),
    .A3(_11839_),
    .ZN(_11917_));
 BUF_X4 _17813_ (.A(_11487_),
    .Z(_11918_));
 AOI211_X2 _17814_ (.A(_11854_),
    .B(_11917_),
    .C1(_11858_),
    .C2(_11918_),
    .ZN(_11919_));
 NOR2_X1 _17815_ (.A1(_11916_),
    .A2(_11919_),
    .ZN(_11920_));
 XNOR2_X2 _17816_ (.A(_11920_),
    .B(_11902_),
    .ZN(\alu_adder_result_ex[10] ));
 CLKBUF_X3 _17817_ (.A(_10673_),
    .Z(_11921_));
 BUF_X4 _17818_ (.A(_11921_),
    .Z(_11922_));
 NOR3_X2 _17819_ (.A1(_10510_),
    .A2(_10374_),
    .A3(net18),
    .ZN(_11923_));
 OAI21_X2 _17820_ (.A(_10386_),
    .B1(_11320_),
    .B2(_11923_),
    .ZN(_11924_));
 NAND2_X4 _17821_ (.A1(_10317_),
    .A2(_11924_),
    .ZN(_11925_));
 MUX2_X2 _17822_ (.A(_11073_),
    .B(_10928_),
    .S(_10926_),
    .Z(_11926_));
 NOR3_X1 _17823_ (.A1(_10346_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_11927_));
 BUF_X8 _17824_ (.A(_10709_),
    .Z(_11928_));
 BUF_X8 _17825_ (.A(_11928_),
    .Z(_11929_));
 BUF_X4 _17826_ (.A(_10432_),
    .Z(_11930_));
 BUF_X4 _17827_ (.A(_10421_),
    .Z(_11931_));
 BUF_X4 _17828_ (.A(_11931_),
    .Z(_11932_));
 BUF_X8 _17829_ (.A(_10466_),
    .Z(_11933_));
 BUF_X8 _17830_ (.A(_11933_),
    .Z(_11934_));
 BUF_X8 _17831_ (.A(_11934_),
    .Z(_11935_));
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 BUF_X32 _17833_ (.A(_10459_),
    .Z(_11937_));
 BUF_X32 _17834_ (.A(_11937_),
    .Z(_11938_));
 BUF_X4 _17835_ (.A(_11938_),
    .Z(_11939_));
 MUX2_X1 _17836_ (.A(_00224_),
    .B(_00226_),
    .S(_11939_),
    .Z(_11940_));
 NOR2_X1 _17837_ (.A1(_11935_),
    .A2(_11940_),
    .ZN(_11941_));
 BUF_X4 _17838_ (.A(_10697_),
    .Z(_11942_));
 BUF_X8 _17839_ (.A(_10459_),
    .Z(_11943_));
 BUF_X4 _17840_ (.A(_11943_),
    .Z(_11944_));
 MUX2_X1 _17841_ (.A(_00225_),
    .B(_00227_),
    .S(_11944_),
    .Z(_11945_));
 NOR2_X1 _17842_ (.A1(_11942_),
    .A2(_11945_),
    .ZN(_11946_));
 NOR3_X1 _17843_ (.A1(_11932_),
    .A2(_11941_),
    .A3(_11946_),
    .ZN(_11947_));
 BUF_X4 _17844_ (.A(_10468_),
    .Z(_11948_));
 BUF_X4 _17845_ (.A(_10964_),
    .Z(_11949_));
 NOR2_X1 _17846_ (.A1(_11944_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .ZN(_11950_));
 BUF_X32 _17847_ (.A(_10459_),
    .Z(_11951_));
 BUF_X4 _17848_ (.A(_11951_),
    .Z(_11952_));
 BUF_X4 _17849_ (.A(_11952_),
    .Z(_11953_));
 AOI21_X1 _17850_ (.A(_11950_),
    .B1(_00219_),
    .B2(_11953_),
    .ZN(_11954_));
 BUF_X4 _17851_ (.A(_10466_),
    .Z(_11955_));
 BUF_X4 _17852_ (.A(_11955_),
    .Z(_11956_));
 AOI221_X2 _17853_ (.A(_11948_),
    .B1(_10820_),
    .B2(_11949_),
    .C1(_11954_),
    .C2(_11956_),
    .ZN(_11957_));
 NOR3_X2 _17854_ (.A1(_11930_),
    .A2(_11947_),
    .A3(_11957_),
    .ZN(_11958_));
 BUF_X4 _17855_ (.A(_10436_),
    .Z(_11959_));
 BUF_X4 _17856_ (.A(net393),
    .Z(_11960_));
 MUX2_X1 _17857_ (.A(_00228_),
    .B(_00230_),
    .S(_11960_),
    .Z(_11961_));
 BUF_X8 _17858_ (.A(_10459_),
    .Z(_11962_));
 MUX2_X1 _17859_ (.A(_00229_),
    .B(_00231_),
    .S(_11962_),
    .Z(_11963_));
 BUF_X4 _17860_ (.A(_10466_),
    .Z(_11964_));
 MUX2_X1 _17861_ (.A(_11961_),
    .B(_11963_),
    .S(_11964_),
    .Z(_11965_));
 MUX2_X1 _17862_ (.A(_00220_),
    .B(_00222_),
    .S(_11962_),
    .Z(_11966_));
 MUX2_X1 _17863_ (.A(_00221_),
    .B(_00223_),
    .S(_11962_),
    .Z(_11967_));
 MUX2_X1 _17864_ (.A(_11966_),
    .B(_11967_),
    .S(_11964_),
    .Z(_11968_));
 BUF_X4 _17865_ (.A(_11931_),
    .Z(_11969_));
 MUX2_X1 _17866_ (.A(_11965_),
    .B(_11968_),
    .S(_11969_),
    .Z(_11970_));
 NOR2_X1 _17867_ (.A1(_11959_),
    .A2(_11970_),
    .ZN(_11971_));
 NOR3_X2 _17868_ (.A1(_11929_),
    .A2(_11958_),
    .A3(_11971_),
    .ZN(_11972_));
 MUX2_X1 _17869_ (.A(_00240_),
    .B(_00242_),
    .S(_11952_),
    .Z(_11973_));
 MUX2_X1 _17870_ (.A(_00241_),
    .B(_00243_),
    .S(_11952_),
    .Z(_11974_));
 BUF_X8 _17871_ (.A(_11933_),
    .Z(_11975_));
 MUX2_X1 _17872_ (.A(_11973_),
    .B(_11974_),
    .S(_11975_),
    .Z(_11976_));
 MUX2_X1 _17873_ (.A(_00232_),
    .B(_00234_),
    .S(_11952_),
    .Z(_11977_));
 BUF_X4 _17874_ (.A(_11951_),
    .Z(_11978_));
 MUX2_X1 _17875_ (.A(_00233_),
    .B(_00235_),
    .S(_11978_),
    .Z(_11979_));
 MUX2_X1 _17876_ (.A(_11977_),
    .B(_11979_),
    .S(_11975_),
    .Z(_11980_));
 MUX2_X1 _17877_ (.A(_11976_),
    .B(_11980_),
    .S(_11932_),
    .Z(_11981_));
 MUX2_X1 _17878_ (.A(_00244_),
    .B(_00246_),
    .S(_11952_),
    .Z(_11982_));
 MUX2_X1 _17879_ (.A(_00245_),
    .B(_00247_),
    .S(_11978_),
    .Z(_11983_));
 MUX2_X1 _17880_ (.A(_11982_),
    .B(_11983_),
    .S(_11975_),
    .Z(_11984_));
 MUX2_X1 _17881_ (.A(_00236_),
    .B(_00238_),
    .S(_11978_),
    .Z(_11985_));
 MUX2_X1 _17882_ (.A(_00237_),
    .B(_00239_),
    .S(_11978_),
    .Z(_11986_));
 MUX2_X1 _17883_ (.A(_11985_),
    .B(_11986_),
    .S(_11975_),
    .Z(_11987_));
 MUX2_X1 _17884_ (.A(_11984_),
    .B(_11987_),
    .S(_11932_),
    .Z(_11988_));
 BUF_X8 _17885_ (.A(_10432_),
    .Z(_11989_));
 MUX2_X1 _17886_ (.A(_11981_),
    .B(_11988_),
    .S(_11989_),
    .Z(_11990_));
 BUF_X8 _17887_ (.A(_11928_),
    .Z(_11991_));
 BUF_X8 _17888_ (.A(_11991_),
    .Z(_11992_));
 AOI21_X4 _17889_ (.A(_11972_),
    .B1(_11990_),
    .B2(_11992_),
    .ZN(_11993_));
 CLKBUF_X3 _17890_ (.A(_10317_),
    .Z(_11994_));
 BUF_X4 _17891_ (.A(_11994_),
    .Z(_11995_));
 OAI221_X2 _17892_ (.A(_11922_),
    .B1(_11925_),
    .B2(_11927_),
    .C1(_11995_),
    .C2(_11993_),
    .ZN(_15937_));
 INV_X1 _17893_ (.A(_15937_),
    .ZN(_15933_));
 NOR3_X1 _17894_ (.A1(_10380_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_11996_));
 BUF_X8 _17895_ (.A(_11951_),
    .Z(_11997_));
 MUX2_X1 _17896_ (.A(_00589_),
    .B(_00591_),
    .S(_11997_),
    .Z(_11998_));
 MUX2_X1 _17897_ (.A(_00590_),
    .B(_00592_),
    .S(_11997_),
    .Z(_11999_));
 BUF_X8 _17898_ (.A(_11933_),
    .Z(_12000_));
 MUX2_X1 _17899_ (.A(_11998_),
    .B(_11999_),
    .S(_12000_),
    .Z(_12001_));
 MUX2_X1 _17900_ (.A(_00581_),
    .B(_00583_),
    .S(_11997_),
    .Z(_12002_));
 MUX2_X1 _17901_ (.A(_00582_),
    .B(_00584_),
    .S(_11997_),
    .Z(_12003_));
 MUX2_X1 _17902_ (.A(_12002_),
    .B(_12003_),
    .S(_12000_),
    .Z(_12004_));
 BUF_X4 _17903_ (.A(_11931_),
    .Z(_12005_));
 MUX2_X1 _17904_ (.A(_12001_),
    .B(_12004_),
    .S(_12005_),
    .Z(_12006_));
 NOR2_X1 _17905_ (.A1(_11989_),
    .A2(_12006_),
    .ZN(_12007_));
 BUF_X8 _17906_ (.A(_11937_),
    .Z(_12008_));
 MUX2_X1 _17907_ (.A(_00593_),
    .B(_00595_),
    .S(_12008_),
    .Z(_12009_));
 BUF_X32 _17908_ (.A(_11937_),
    .Z(_12010_));
 MUX2_X1 _17909_ (.A(_00594_),
    .B(_00596_),
    .S(_12010_),
    .Z(_12011_));
 BUF_X4 _17910_ (.A(_11933_),
    .Z(_12012_));
 MUX2_X1 _17911_ (.A(_12009_),
    .B(_12011_),
    .S(_12012_),
    .Z(_12013_));
 MUX2_X1 _17912_ (.A(_00585_),
    .B(_00587_),
    .S(_12010_),
    .Z(_12014_));
 MUX2_X1 _17913_ (.A(_00586_),
    .B(_00588_),
    .S(_12010_),
    .Z(_12015_));
 MUX2_X1 _17914_ (.A(_12014_),
    .B(_12015_),
    .S(_12012_),
    .Z(_12016_));
 BUF_X4 _17915_ (.A(_11931_),
    .Z(_12017_));
 MUX2_X1 _17916_ (.A(_12013_),
    .B(_12016_),
    .S(_12017_),
    .Z(_12018_));
 NOR2_X2 _17917_ (.A1(_11959_),
    .A2(_12018_),
    .ZN(_12019_));
 NOR3_X2 _17918_ (.A1(_10474_),
    .A2(_12007_),
    .A3(_12019_),
    .ZN(_12020_));
 BUF_X8 _17919_ (.A(_11951_),
    .Z(_12021_));
 MUX2_X1 _17920_ (.A(_00577_),
    .B(_00579_),
    .S(_12021_),
    .Z(_12022_));
 BUF_X4 _17921_ (.A(_11951_),
    .Z(_12023_));
 MUX2_X1 _17922_ (.A(_00578_),
    .B(_00580_),
    .S(_12023_),
    .Z(_12024_));
 MUX2_X1 _17923_ (.A(_12022_),
    .B(_12024_),
    .S(_11934_),
    .Z(_12025_));
 MUX2_X1 _17924_ (.A(_00569_),
    .B(_00571_),
    .S(_12023_),
    .Z(_12026_));
 MUX2_X1 _17925_ (.A(_00570_),
    .B(_00572_),
    .S(_12023_),
    .Z(_12027_));
 MUX2_X1 _17926_ (.A(_12026_),
    .B(_12027_),
    .S(_11934_),
    .Z(_12028_));
 BUF_X4 _17927_ (.A(_11931_),
    .Z(_12029_));
 MUX2_X1 _17928_ (.A(_12025_),
    .B(_12028_),
    .S(_12029_),
    .Z(_12030_));
 NOR2_X1 _17929_ (.A1(_11959_),
    .A2(_12030_),
    .ZN(_12031_));
 INV_X1 _17930_ (.A(_00567_),
    .ZN(_12032_));
 NOR2_X1 _17931_ (.A1(_11953_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .ZN(_12033_));
 BUF_X8 _17932_ (.A(_11939_),
    .Z(_12034_));
 AOI21_X1 _17933_ (.A(_12033_),
    .B1(_00568_),
    .B2(_12034_),
    .ZN(_12035_));
 AOI221_X1 _17934_ (.A(_11948_),
    .B1(_12032_),
    .B2(_11949_),
    .C1(_12035_),
    .C2(_11956_),
    .ZN(_12036_));
 BUF_X8 _17935_ (.A(_11944_),
    .Z(_12037_));
 MUX2_X1 _17936_ (.A(_00573_),
    .B(_00575_),
    .S(_12037_),
    .Z(_12038_));
 MUX2_X1 _17937_ (.A(_00574_),
    .B(_00576_),
    .S(_12037_),
    .Z(_12039_));
 MUX2_X1 _17938_ (.A(_12038_),
    .B(_12039_),
    .S(_11935_),
    .Z(_12040_));
 BUF_X8 _17939_ (.A(_11948_),
    .Z(_12041_));
 AOI21_X1 _17940_ (.A(_12036_),
    .B1(_12040_),
    .B2(_12041_),
    .ZN(_12042_));
 AOI21_X2 _17941_ (.A(_12031_),
    .B1(_12042_),
    .B2(_11959_),
    .ZN(_12043_));
 AOI21_X4 _17942_ (.A(_12020_),
    .B1(_12043_),
    .B2(_10474_),
    .ZN(_12044_));
 OAI221_X2 _17943_ (.A(_11922_),
    .B1(_11925_),
    .B2(_11996_),
    .C1(_11995_),
    .C2(_12044_),
    .ZN(_15945_));
 INV_X1 _17944_ (.A(_15945_),
    .ZN(_15941_));
 NAND2_X1 _17945_ (.A1(_10621_),
    .A2(_00568_),
    .ZN(_12045_));
 OAI21_X1 _17946_ (.A(_12045_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .B2(_10602_),
    .ZN(_12046_));
 OAI221_X1 _17947_ (.A(_10570_),
    .B1(_00567_),
    .B2(_10757_),
    .C1(_12046_),
    .C2(_10580_),
    .ZN(_12047_));
 MUX2_X1 _17948_ (.A(_00573_),
    .B(_00575_),
    .S(_11546_),
    .Z(_12048_));
 MUX2_X1 _17949_ (.A(_00574_),
    .B(_00576_),
    .S(_10823_),
    .Z(_12049_));
 MUX2_X1 _17950_ (.A(_12048_),
    .B(_12049_),
    .S(_11535_),
    .Z(_12050_));
 AOI21_X1 _17951_ (.A(_10831_),
    .B1(_12050_),
    .B2(_10766_),
    .ZN(_12051_));
 NAND2_X1 _17952_ (.A1(_12047_),
    .A2(_12051_),
    .ZN(_12052_));
 MUX2_X1 _17953_ (.A(_00589_),
    .B(_00591_),
    .S(_10585_),
    .Z(_12053_));
 MUX2_X1 _17954_ (.A(_00590_),
    .B(_00592_),
    .S(_10585_),
    .Z(_12054_));
 MUX2_X1 _17955_ (.A(_12053_),
    .B(_12054_),
    .S(_10787_),
    .Z(_12055_));
 MUX2_X1 _17956_ (.A(_00581_),
    .B(_00583_),
    .S(_10619_),
    .Z(_12056_));
 MUX2_X1 _17957_ (.A(_00582_),
    .B(_00584_),
    .S(_10619_),
    .Z(_12057_));
 MUX2_X1 _17958_ (.A(_12056_),
    .B(_12057_),
    .S(_10787_),
    .Z(_12058_));
 MUX2_X1 _17959_ (.A(_12055_),
    .B(_12058_),
    .S(_10828_),
    .Z(_12059_));
 MUX2_X1 _17960_ (.A(_00593_),
    .B(_00595_),
    .S(_11639_),
    .Z(_12060_));
 MUX2_X1 _17961_ (.A(_00594_),
    .B(_00596_),
    .S(_11678_),
    .Z(_12061_));
 MUX2_X1 _17962_ (.A(_12060_),
    .B(_12061_),
    .S(_10626_),
    .Z(_12062_));
 MUX2_X1 _17963_ (.A(_00585_),
    .B(_00587_),
    .S(_11678_),
    .Z(_12063_));
 MUX2_X1 _17964_ (.A(_00586_),
    .B(_00588_),
    .S(_11678_),
    .Z(_12064_));
 MUX2_X1 _17965_ (.A(_12063_),
    .B(_12064_),
    .S(_10626_),
    .Z(_12065_));
 MUX2_X1 _17966_ (.A(_12062_),
    .B(_12065_),
    .S(_10827_),
    .Z(_12066_));
 MUX2_X1 _17967_ (.A(_00577_),
    .B(_00579_),
    .S(_11678_),
    .Z(_12067_));
 MUX2_X1 _17968_ (.A(_00578_),
    .B(_00580_),
    .S(_11678_),
    .Z(_12068_));
 MUX2_X1 _17969_ (.A(_12067_),
    .B(_12068_),
    .S(_10626_),
    .Z(_12069_));
 MUX2_X1 _17970_ (.A(_00569_),
    .B(_00571_),
    .S(_11678_),
    .Z(_12070_));
 MUX2_X1 _17971_ (.A(_00570_),
    .B(_00572_),
    .S(_11678_),
    .Z(_12071_));
 MUX2_X1 _17972_ (.A(_12070_),
    .B(_12071_),
    .S(_10786_),
    .Z(_12072_));
 MUX2_X1 _17973_ (.A(_12069_),
    .B(_12072_),
    .S(_10827_),
    .Z(_12073_));
 MUX2_X1 _17974_ (.A(_12066_),
    .B(_12073_),
    .S(_10574_),
    .Z(_12074_));
 OAI221_X2 _17975_ (.A(_12052_),
    .B1(_12059_),
    .B2(_11371_),
    .C1(_12074_),
    .C2(_10609_),
    .ZN(_12075_));
 BUF_X1 _17976_ (.A(\cs_registers_i.pc_id_i[13] ),
    .Z(_12076_));
 AND2_X1 _17977_ (.A1(_12076_),
    .A2(_11593_),
    .ZN(_12077_));
 AOI222_X2 _17978_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(_10397_),
    .B1(_10816_),
    .B2(_12075_),
    .C1(_12077_),
    .C2(_10870_),
    .ZN(_12078_));
 BUF_X4 _17979_ (.A(_12078_),
    .Z(_15944_));
 CLKBUF_X2 _17980_ (.A(_15422_),
    .Z(_12079_));
 INV_X2 _17981_ (.A(_12079_),
    .ZN(_12080_));
 INV_X1 _17982_ (.A(_15417_),
    .ZN(_12081_));
 BUF_X1 rebuffer42 (.A(_13155_),
    .Z(net313));
 BUF_X1 _17984_ (.A(_15413_),
    .Z(_12083_));
 OAI21_X1 _17985_ (.A(_15418_),
    .B1(_12083_),
    .B2(_11910_),
    .ZN(_12084_));
 NAND2_X1 _17986_ (.A1(_12081_),
    .A2(_12084_),
    .ZN(_12085_));
 XNOR2_X2 _17987_ (.A(_12080_),
    .B(_12085_),
    .ZN(\alu_adder_result_ex[13] ));
 NAND2_X1 _17988_ (.A1(_11902_),
    .A2(_11900_),
    .ZN(_12086_));
 NOR2_X2 _17989_ (.A1(_11905_),
    .A2(_12086_),
    .ZN(_12087_));
 NAND3_X1 _17990_ (.A1(net368),
    .A2(_11860_),
    .A3(_12087_),
    .ZN(_12088_));
 OAI21_X1 _17991_ (.A(_11908_),
    .B1(_11904_),
    .B2(_11903_),
    .ZN(_12089_));
 AND2_X1 _17992_ (.A1(_11900_),
    .A2(_12089_),
    .ZN(_12090_));
 OR2_X1 _17993_ (.A1(_12083_),
    .A2(_12090_),
    .ZN(_12091_));
 OR3_X1 _17994_ (.A1(net367),
    .A2(_11839_),
    .A3(_12091_),
    .ZN(_12092_));
 NAND3_X1 _17995_ (.A1(net367),
    .A2(_11839_),
    .A3(_12087_),
    .ZN(_12093_));
 OAI221_X2 _17996_ (.A(_12088_),
    .B1(_12092_),
    .B2(_11860_),
    .C1(_12093_),
    .C2(_11863_),
    .ZN(_12094_));
 NOR3_X1 _17997_ (.A1(net368),
    .A2(_12091_),
    .A3(_12087_),
    .ZN(_12095_));
 INV_X1 _17998_ (.A(net449),
    .ZN(_12096_));
 NOR2_X1 _17999_ (.A1(_12083_),
    .A2(_12090_),
    .ZN(_12097_));
 NOR2_X1 _18000_ (.A1(_12096_),
    .A2(_12097_),
    .ZN(_12098_));
 AOI21_X4 _18001_ (.A(_11854_),
    .B1(_11918_),
    .B2(_11858_),
    .ZN(_12099_));
 NOR4_X2 _18002_ (.A1(net367),
    .A2(_12099_),
    .A3(_11860_),
    .A4(_12091_),
    .ZN(_12100_));
 NOR4_X2 _18003_ (.A1(_12094_),
    .A2(_12095_),
    .A3(_12098_),
    .A4(_12100_),
    .ZN(_12101_));
 BUF_X4 _18004_ (.A(_12101_),
    .Z(\alu_adder_result_ex[12] ));
 BUF_X4 _18005_ (.A(_11432_),
    .Z(_12102_));
 BUF_X4 _18006_ (.A(_12102_),
    .Z(_12103_));
 NOR3_X1 _18007_ (.A1(_12103_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12104_));
 MUX2_X1 _18008_ (.A(_00604_),
    .B(_00606_),
    .S(_11944_),
    .Z(_12105_));
 NOR2_X1 _18009_ (.A1(_11956_),
    .A2(_12105_),
    .ZN(_12106_));
 MUX2_X1 _18010_ (.A(_00605_),
    .B(_00607_),
    .S(_11944_),
    .Z(_12107_));
 NOR2_X1 _18011_ (.A1(_11942_),
    .A2(_12107_),
    .ZN(_12108_));
 NOR3_X1 _18012_ (.A1(_11932_),
    .A2(_12106_),
    .A3(_12108_),
    .ZN(_12109_));
 INV_X1 _18013_ (.A(_00598_),
    .ZN(_12110_));
 BUF_X4 _18014_ (.A(net393),
    .Z(_12111_));
 BUF_X4 _18015_ (.A(_12111_),
    .Z(_12112_));
 NOR2_X1 _18016_ (.A1(_12112_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .ZN(_12113_));
 AOI21_X1 _18017_ (.A(_12113_),
    .B1(_00599_),
    .B2(_11939_),
    .ZN(_12114_));
 AOI221_X2 _18018_ (.A(_10468_),
    .B1(_12110_),
    .B2(_11949_),
    .C1(_12114_),
    .C2(_11975_),
    .ZN(_12115_));
 NOR3_X1 _18019_ (.A1(_11930_),
    .A2(_12109_),
    .A3(_12115_),
    .ZN(_12116_));
 BUF_X4 _18020_ (.A(_10436_),
    .Z(_12117_));
 MUX2_X1 _18021_ (.A(_00608_),
    .B(_00610_),
    .S(_11943_),
    .Z(_12118_));
 MUX2_X1 _18022_ (.A(_00609_),
    .B(_00611_),
    .S(_11943_),
    .Z(_12119_));
 MUX2_X1 _18023_ (.A(_12118_),
    .B(_12119_),
    .S(_11955_),
    .Z(_12120_));
 MUX2_X1 _18024_ (.A(_00600_),
    .B(_00602_),
    .S(_11943_),
    .Z(_12121_));
 MUX2_X1 _18025_ (.A(_00601_),
    .B(_00603_),
    .S(_11943_),
    .Z(_12122_));
 MUX2_X1 _18026_ (.A(_12121_),
    .B(_12122_),
    .S(_11955_),
    .Z(_12123_));
 BUF_X4 _18027_ (.A(_11931_),
    .Z(_12124_));
 MUX2_X1 _18028_ (.A(_12120_),
    .B(_12123_),
    .S(_12124_),
    .Z(_12125_));
 NOR2_X1 _18029_ (.A1(_12117_),
    .A2(_12125_),
    .ZN(_12126_));
 NOR3_X2 _18030_ (.A1(_11991_),
    .A2(_12116_),
    .A3(_12126_),
    .ZN(_12127_));
 MUX2_X1 _18031_ (.A(_00620_),
    .B(_00622_),
    .S(_11997_),
    .Z(_12128_));
 BUF_X8 _18032_ (.A(_11951_),
    .Z(_12129_));
 MUX2_X1 _18033_ (.A(_00621_),
    .B(_00623_),
    .S(_12129_),
    .Z(_12130_));
 MUX2_X1 _18034_ (.A(_12128_),
    .B(_12130_),
    .S(_12000_),
    .Z(_12131_));
 MUX2_X1 _18035_ (.A(_00612_),
    .B(_00614_),
    .S(_11997_),
    .Z(_12132_));
 MUX2_X1 _18036_ (.A(_00613_),
    .B(_00615_),
    .S(_12129_),
    .Z(_12133_));
 MUX2_X1 _18037_ (.A(_12132_),
    .B(_12133_),
    .S(_12000_),
    .Z(_12134_));
 MUX2_X1 _18038_ (.A(_12131_),
    .B(_12134_),
    .S(_12005_),
    .Z(_12135_));
 MUX2_X1 _18039_ (.A(_00624_),
    .B(_00626_),
    .S(_12129_),
    .Z(_12136_));
 MUX2_X1 _18040_ (.A(_00625_),
    .B(_00627_),
    .S(_12129_),
    .Z(_12137_));
 MUX2_X1 _18041_ (.A(_12136_),
    .B(_12137_),
    .S(_12000_),
    .Z(_12138_));
 MUX2_X1 _18042_ (.A(_00616_),
    .B(_00618_),
    .S(_12129_),
    .Z(_12139_));
 MUX2_X1 _18043_ (.A(_00617_),
    .B(_00619_),
    .S(_12129_),
    .Z(_12140_));
 MUX2_X1 _18044_ (.A(_12139_),
    .B(_12140_),
    .S(_12000_),
    .Z(_12141_));
 MUX2_X1 _18045_ (.A(_12138_),
    .B(_12141_),
    .S(_12005_),
    .Z(_12142_));
 MUX2_X1 _18046_ (.A(_12135_),
    .B(_12142_),
    .S(_11930_),
    .Z(_12143_));
 AOI21_X4 _18047_ (.A(_12127_),
    .B1(_12143_),
    .B2(_11992_),
    .ZN(_12144_));
 OAI221_X2 _18048_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12104_),
    .C1(_12144_),
    .C2(_11995_),
    .ZN(_15953_));
 INV_X1 _18049_ (.A(_15953_),
    .ZN(_15949_));
 MUX2_X1 _18050_ (.A(_00604_),
    .B(_00606_),
    .S(_11363_),
    .Z(_12145_));
 MUX2_X1 _18051_ (.A(_00605_),
    .B(_00607_),
    .S(_11363_),
    .Z(_12146_));
 MUX2_X1 _18052_ (.A(_12145_),
    .B(_12146_),
    .S(_11366_),
    .Z(_12147_));
 NOR2_X1 _18053_ (.A1(_10620_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .ZN(_12148_));
 AOI21_X1 _18054_ (.A(_12148_),
    .B1(_00599_),
    .B2(_10601_),
    .ZN(_12149_));
 AOI22_X1 _18055_ (.A1(_12110_),
    .A2(_10822_),
    .B1(_12149_),
    .B2(_10788_),
    .ZN(_12150_));
 MUX2_X1 _18056_ (.A(_12147_),
    .B(_12150_),
    .S(_11358_),
    .Z(_12151_));
 MUX2_X1 _18057_ (.A(_00616_),
    .B(_00618_),
    .S(_11546_),
    .Z(_12152_));
 MUX2_X1 _18058_ (.A(_00617_),
    .B(_00619_),
    .S(_11546_),
    .Z(_12153_));
 MUX2_X1 _18059_ (.A(_12152_),
    .B(_12153_),
    .S(_10595_),
    .Z(_12154_));
 NAND2_X1 _18060_ (.A1(_10778_),
    .A2(_12154_),
    .ZN(_12155_));
 MUX2_X1 _18061_ (.A(_00614_),
    .B(_00615_),
    .S(_10595_),
    .Z(_12156_));
 NAND2_X1 _18062_ (.A1(_10794_),
    .A2(_12156_),
    .ZN(_12157_));
 MUX2_X1 _18063_ (.A(_00612_),
    .B(_00613_),
    .S(_11877_),
    .Z(_12158_));
 AOI21_X1 _18064_ (.A(_10575_),
    .B1(_10785_),
    .B2(_12158_),
    .ZN(_12159_));
 NAND3_X1 _18065_ (.A1(_12155_),
    .A2(_12157_),
    .A3(_12159_),
    .ZN(_12160_));
 MUX2_X1 _18066_ (.A(_00620_),
    .B(_00621_),
    .S(_10787_),
    .Z(_12161_));
 NOR3_X1 _18067_ (.A1(_10622_),
    .A2(_11676_),
    .A3(_12161_),
    .ZN(_12162_));
 MUX2_X1 _18068_ (.A(_00622_),
    .B(_00623_),
    .S(_11534_),
    .Z(_12163_));
 NOR3_X1 _18069_ (.A1(_10632_),
    .A2(_10751_),
    .A3(_12163_),
    .ZN(_12164_));
 MUX2_X1 _18070_ (.A(_00624_),
    .B(_00625_),
    .S(_10593_),
    .Z(_12165_));
 MUX2_X1 _18071_ (.A(_00626_),
    .B(_00627_),
    .S(_10593_),
    .Z(_12166_));
 MUX2_X1 _18072_ (.A(_12165_),
    .B(_12166_),
    .S(_10614_),
    .Z(_12167_));
 OAI21_X1 _18073_ (.A(_10765_),
    .B1(_12167_),
    .B2(_11775_),
    .ZN(_12168_));
 NOR3_X1 _18074_ (.A1(_12162_),
    .A2(_12164_),
    .A3(_12168_),
    .ZN(_12169_));
 MUX2_X1 _18075_ (.A(_00608_),
    .B(_00610_),
    .S(_10613_),
    .Z(_12170_));
 MUX2_X1 _18076_ (.A(_00609_),
    .B(_00611_),
    .S(_10613_),
    .Z(_12171_));
 MUX2_X1 _18077_ (.A(_12170_),
    .B(_12171_),
    .S(_10796_),
    .Z(_12172_));
 MUX2_X1 _18078_ (.A(_00600_),
    .B(_00602_),
    .S(_10613_),
    .Z(_12173_));
 MUX2_X1 _18079_ (.A(_00601_),
    .B(_00603_),
    .S(_10613_),
    .Z(_12174_));
 MUX2_X1 _18080_ (.A(_12173_),
    .B(_12174_),
    .S(_10796_),
    .Z(_12175_));
 MUX2_X1 _18081_ (.A(_12172_),
    .B(_12175_),
    .S(_10828_),
    .Z(_12176_));
 OAI222_X2 _18082_ (.A1(_10831_),
    .A2(_12151_),
    .B1(_12160_),
    .B2(_12169_),
    .C1(_12176_),
    .C2(_10855_),
    .ZN(_12177_));
 NAND2_X1 _18083_ (.A1(_11596_),
    .A2(_12177_),
    .ZN(_12178_));
 CLKBUF_X2 _18084_ (.A(\cs_registers_i.pc_id_i[14] ),
    .Z(_12179_));
 AND2_X1 _18085_ (.A1(_12179_),
    .A2(_11593_),
    .ZN(_12180_));
 AOI22_X2 _18086_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(_10741_),
    .B1(_10870_),
    .B2(_12180_),
    .ZN(_12181_));
 NAND2_X1 _18087_ (.A1(_12178_),
    .A2(_12181_),
    .ZN(_15948_));
 INV_X2 _18088_ (.A(_15948_),
    .ZN(_15952_));
 NOR3_X1 _18089_ (.A1(_10582_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12182_));
 MUX2_X1 _18090_ (.A(_00635_),
    .B(_00637_),
    .S(_11944_),
    .Z(_12183_));
 NOR2_X1 _18091_ (.A1(_11935_),
    .A2(_12183_),
    .ZN(_12184_));
 MUX2_X1 _18092_ (.A(_00636_),
    .B(_00638_),
    .S(_11944_),
    .Z(_12185_));
 NOR2_X1 _18093_ (.A1(_11942_),
    .A2(_12185_),
    .ZN(_12186_));
 NOR3_X1 _18094_ (.A1(_11932_),
    .A2(_12184_),
    .A3(_12186_),
    .ZN(_12187_));
 INV_X1 _18095_ (.A(_00629_),
    .ZN(_12188_));
 NOR2_X1 _18096_ (.A1(_11944_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .ZN(_12189_));
 AOI21_X1 _18097_ (.A(_12189_),
    .B1(_00630_),
    .B2(_11953_),
    .ZN(_12190_));
 AOI221_X1 _18098_ (.A(_11948_),
    .B1(_12188_),
    .B2(_11949_),
    .C1(_12190_),
    .C2(_11975_),
    .ZN(_12191_));
 NOR3_X1 _18099_ (.A1(_11930_),
    .A2(_12187_),
    .A3(_12191_),
    .ZN(_12192_));
 MUX2_X1 _18100_ (.A(_00639_),
    .B(_00641_),
    .S(_11943_),
    .Z(_12193_));
 BUF_X4 _18101_ (.A(net393),
    .Z(_12194_));
 MUX2_X1 _18102_ (.A(_00640_),
    .B(_00642_),
    .S(_12194_),
    .Z(_12195_));
 MUX2_X1 _18103_ (.A(_12193_),
    .B(_12195_),
    .S(_11955_),
    .Z(_12196_));
 MUX2_X1 _18104_ (.A(_00631_),
    .B(_00633_),
    .S(_12194_),
    .Z(_12197_));
 MUX2_X1 _18105_ (.A(_00632_),
    .B(_00634_),
    .S(_12194_),
    .Z(_12198_));
 MUX2_X1 _18106_ (.A(_12197_),
    .B(_12198_),
    .S(_11955_),
    .Z(_12199_));
 BUF_X4 _18107_ (.A(_11931_),
    .Z(_12200_));
 MUX2_X1 _18108_ (.A(_12196_),
    .B(_12199_),
    .S(_12200_),
    .Z(_12201_));
 NOR2_X1 _18109_ (.A1(_12117_),
    .A2(_12201_),
    .ZN(_12202_));
 NOR3_X2 _18110_ (.A1(_11991_),
    .A2(_12192_),
    .A3(_12202_),
    .ZN(_12203_));
 BUF_X8 _18111_ (.A(_11951_),
    .Z(_12204_));
 MUX2_X1 _18112_ (.A(_00651_),
    .B(_00653_),
    .S(_12204_),
    .Z(_12205_));
 MUX2_X1 _18113_ (.A(_00652_),
    .B(_00654_),
    .S(_12204_),
    .Z(_12206_));
 BUF_X16 _18114_ (.A(_11933_),
    .Z(_12207_));
 MUX2_X1 _18115_ (.A(_12205_),
    .B(_12206_),
    .S(_12207_),
    .Z(_12208_));
 MUX2_X1 _18116_ (.A(_00643_),
    .B(_00645_),
    .S(_12204_),
    .Z(_12209_));
 MUX2_X1 _18117_ (.A(_00644_),
    .B(_00646_),
    .S(_12021_),
    .Z(_12210_));
 MUX2_X1 _18118_ (.A(_12209_),
    .B(_12210_),
    .S(_11934_),
    .Z(_12211_));
 MUX2_X1 _18119_ (.A(_12208_),
    .B(_12211_),
    .S(_12029_),
    .Z(_12212_));
 MUX2_X1 _18120_ (.A(_00655_),
    .B(_00657_),
    .S(_12021_),
    .Z(_12213_));
 MUX2_X1 _18121_ (.A(_00656_),
    .B(_00658_),
    .S(_12021_),
    .Z(_12214_));
 MUX2_X1 _18122_ (.A(_12213_),
    .B(_12214_),
    .S(_11934_),
    .Z(_12215_));
 MUX2_X1 _18123_ (.A(_00647_),
    .B(_00649_),
    .S(_12021_),
    .Z(_12216_));
 MUX2_X1 _18124_ (.A(_00648_),
    .B(_00650_),
    .S(_12021_),
    .Z(_12217_));
 MUX2_X1 _18125_ (.A(_12216_),
    .B(_12217_),
    .S(_11934_),
    .Z(_12218_));
 MUX2_X1 _18126_ (.A(_12215_),
    .B(_12218_),
    .S(_12029_),
    .Z(_12219_));
 MUX2_X1 _18127_ (.A(_12212_),
    .B(_12219_),
    .S(_11989_),
    .Z(_12220_));
 AOI21_X4 _18128_ (.A(_12203_),
    .B1(_11992_),
    .B2(_12220_),
    .ZN(_12221_));
 OAI221_X2 _18129_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12182_),
    .C1(_12221_),
    .C2(_11995_),
    .ZN(_15956_));
 INV_X1 _18130_ (.A(_15956_),
    .ZN(_15960_));
 MUX2_X1 _18131_ (.A(_00655_),
    .B(_00657_),
    .S(_11372_),
    .Z(_12222_));
 MUX2_X1 _18132_ (.A(_00656_),
    .B(_00658_),
    .S(_10599_),
    .Z(_12223_));
 MUX2_X1 _18133_ (.A(_12222_),
    .B(_12223_),
    .S(_11375_),
    .Z(_12224_));
 MUX2_X1 _18134_ (.A(_00647_),
    .B(_00649_),
    .S(_10599_),
    .Z(_12225_));
 MUX2_X1 _18135_ (.A(_00648_),
    .B(_00650_),
    .S(_10599_),
    .Z(_12226_));
 MUX2_X1 _18136_ (.A(_12225_),
    .B(_12226_),
    .S(_11375_),
    .Z(_12227_));
 MUX2_X1 _18137_ (.A(_12224_),
    .B(_12227_),
    .S(_10569_),
    .Z(_12228_));
 MUX2_X1 _18138_ (.A(_00651_),
    .B(_00653_),
    .S(_10599_),
    .Z(_12229_));
 MUX2_X1 _18139_ (.A(_00652_),
    .B(_00654_),
    .S(_10599_),
    .Z(_12230_));
 MUX2_X1 _18140_ (.A(_12229_),
    .B(_12230_),
    .S(_11375_),
    .Z(_12231_));
 MUX2_X1 _18141_ (.A(_00643_),
    .B(_00645_),
    .S(_10599_),
    .Z(_12232_));
 MUX2_X1 _18142_ (.A(_00644_),
    .B(_00646_),
    .S(_10599_),
    .Z(_12233_));
 MUX2_X1 _18143_ (.A(_12232_),
    .B(_12233_),
    .S(_11534_),
    .Z(_12234_));
 MUX2_X1 _18144_ (.A(_12231_),
    .B(_12234_),
    .S(_10569_),
    .Z(_12235_));
 MUX2_X1 _18145_ (.A(_12228_),
    .B(_12235_),
    .S(_10608_),
    .Z(_12236_));
 MUX2_X1 _18146_ (.A(_00639_),
    .B(_00641_),
    .S(_10620_),
    .Z(_12237_));
 MUX2_X1 _18147_ (.A(_00640_),
    .B(_00642_),
    .S(_10620_),
    .Z(_12238_));
 MUX2_X1 _18148_ (.A(_12237_),
    .B(_12238_),
    .S(_10788_),
    .Z(_12239_));
 NAND2_X1 _18149_ (.A1(_11533_),
    .A2(_12239_),
    .ZN(_12240_));
 MUX2_X1 _18150_ (.A(_00631_),
    .B(_00633_),
    .S(_10620_),
    .Z(_12241_));
 MUX2_X1 _18151_ (.A(_00632_),
    .B(_00634_),
    .S(_10620_),
    .Z(_12242_));
 MUX2_X1 _18152_ (.A(_12241_),
    .B(_12242_),
    .S(_10788_),
    .Z(_12243_));
 NAND2_X1 _18153_ (.A1(_10570_),
    .A2(_12243_),
    .ZN(_12244_));
 NAND3_X2 _18154_ (.A1(_10752_),
    .A2(_12240_),
    .A3(_12244_),
    .ZN(_12245_));
 NAND2_X1 _18155_ (.A1(_10615_),
    .A2(_00630_),
    .ZN(_12246_));
 OAI21_X1 _18156_ (.A(_12246_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B2(_10589_),
    .ZN(_12247_));
 OAI221_X2 _18157_ (.A(_10570_),
    .B1(_00629_),
    .B2(_10757_),
    .C1(_12247_),
    .C2(_10581_),
    .ZN(_12248_));
 MUX2_X1 _18158_ (.A(_00635_),
    .B(_00637_),
    .S(_10823_),
    .Z(_12249_));
 MUX2_X1 _18159_ (.A(_00636_),
    .B(_00638_),
    .S(_10600_),
    .Z(_12250_));
 MUX2_X1 _18160_ (.A(_12249_),
    .B(_12250_),
    .S(_11535_),
    .Z(_12251_));
 AOI21_X1 _18161_ (.A(_11676_),
    .B1(_10766_),
    .B2(_12251_),
    .ZN(_12252_));
 AOI21_X2 _18162_ (.A(_10749_),
    .B1(_12248_),
    .B2(_12252_),
    .ZN(_12253_));
 AOI22_X4 _18163_ (.A1(_10750_),
    .A2(_12236_),
    .B1(_12245_),
    .B2(_12253_),
    .ZN(_12254_));
 NAND2_X1 _18164_ (.A1(_11596_),
    .A2(_12254_),
    .ZN(_12255_));
 AND2_X1 _18165_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_11593_),
    .ZN(_12256_));
 AOI22_X4 _18166_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(_10741_),
    .B1(_10683_),
    .B2(_12256_),
    .ZN(_12257_));
 NAND2_X4 _18167_ (.A1(_12255_),
    .A2(_12257_),
    .ZN(_15961_));
 INV_X2 _18168_ (.A(_15961_),
    .ZN(_15957_));
 INV_X1 _18169_ (.A(_15430_),
    .ZN(_12258_));
 INV_X1 _18170_ (.A(_15421_),
    .ZN(_12259_));
 AOI21_X2 _18171_ (.A(_15417_),
    .B1(_12083_),
    .B2(_15418_),
    .ZN(_12260_));
 OAI21_X2 _18172_ (.A(_12259_),
    .B1(_12260_),
    .B2(_12080_),
    .ZN(_12261_));
 BUF_X2 _18173_ (.A(_15426_),
    .Z(_12262_));
 AOI21_X2 _18174_ (.A(_15425_),
    .B1(_12261_),
    .B2(_12262_),
    .ZN(_12263_));
 NAND3_X1 _18175_ (.A1(net449),
    .A2(_12079_),
    .A3(_12262_),
    .ZN(_12264_));
 NAND3_X1 _18176_ (.A1(_12258_),
    .A2(_12263_),
    .A3(_12264_),
    .ZN(_12265_));
 OAI21_X2 _18177_ (.A(_12265_),
    .B1(_12263_),
    .B2(_12258_),
    .ZN(_12266_));
 NAND2_X2 _18178_ (.A1(net449),
    .A2(_12079_),
    .ZN(_12267_));
 NAND2_X2 _18179_ (.A1(_12262_),
    .A2(_15430_),
    .ZN(_12268_));
 NOR2_X2 _18180_ (.A1(_12267_),
    .A2(_12268_),
    .ZN(_12269_));
 AND2_X1 _18181_ (.A1(_11910_),
    .A2(_12269_),
    .ZN(_12270_));
 NAND2_X1 _18182_ (.A1(_12258_),
    .A2(_12263_),
    .ZN(_12271_));
 NOR2_X1 _18183_ (.A1(_11910_),
    .A2(_12271_),
    .ZN(_12272_));
 OR2_X2 _18184_ (.A1(_12270_),
    .A2(_12272_),
    .ZN(_12273_));
 NOR2_X4 _18185_ (.A1(_12266_),
    .A2(_12273_),
    .ZN(\alu_adder_result_ex[15] ));
 AOI21_X1 _18186_ (.A(_12083_),
    .B1(_11901_),
    .B2(_11900_),
    .ZN(_12274_));
 OAI21_X1 _18187_ (.A(_12081_),
    .B1(_12274_),
    .B2(_12096_),
    .ZN(_12275_));
 AOI21_X1 _18188_ (.A(_15421_),
    .B1(_12275_),
    .B2(_12079_),
    .ZN(_12276_));
 OAI21_X1 _18189_ (.A(_12276_),
    .B1(_12267_),
    .B2(_12086_),
    .ZN(_12277_));
 INV_X1 _18190_ (.A(_12276_),
    .ZN(_12278_));
 OR2_X1 _18191_ (.A1(_11916_),
    .A2(_12278_),
    .ZN(_12279_));
 OAI21_X2 _18192_ (.A(_12277_),
    .B1(_12279_),
    .B2(_11919_),
    .ZN(_12280_));
 XNOR2_X2 _18193_ (.A(_12280_),
    .B(_12262_),
    .ZN(\alu_adder_result_ex[14] ));
 NOR3_X1 _18194_ (.A1(_10632_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12281_));
 MUX2_X1 _18195_ (.A(_00666_),
    .B(_00668_),
    .S(_11944_),
    .Z(_12282_));
 NOR2_X1 _18196_ (.A1(_11935_),
    .A2(_12282_),
    .ZN(_12283_));
 MUX2_X1 _18197_ (.A(_00667_),
    .B(_00669_),
    .S(_11944_),
    .Z(_12284_));
 NOR2_X1 _18198_ (.A1(_11942_),
    .A2(_12284_),
    .ZN(_12285_));
 NOR3_X1 _18199_ (.A1(_11932_),
    .A2(_12283_),
    .A3(_12285_),
    .ZN(_12286_));
 INV_X1 _18200_ (.A(_00660_),
    .ZN(_12287_));
 NOR2_X1 _18201_ (.A1(_12112_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .ZN(_12288_));
 AOI21_X1 _18202_ (.A(_12288_),
    .B1(_00661_),
    .B2(_11953_),
    .ZN(_12289_));
 AOI221_X1 _18203_ (.A(_11948_),
    .B1(_12287_),
    .B2(_11949_),
    .C1(_12289_),
    .C2(_11975_),
    .ZN(_12290_));
 NOR3_X1 _18204_ (.A1(_11930_),
    .A2(_12286_),
    .A3(_12290_),
    .ZN(_12291_));
 MUX2_X1 _18205_ (.A(_00670_),
    .B(_00672_),
    .S(_11943_),
    .Z(_12292_));
 MUX2_X1 _18206_ (.A(_00671_),
    .B(_00673_),
    .S(_11943_),
    .Z(_12293_));
 MUX2_X1 _18207_ (.A(_12292_),
    .B(_12293_),
    .S(_11955_),
    .Z(_12294_));
 MUX2_X1 _18208_ (.A(_00662_),
    .B(_00664_),
    .S(_12194_),
    .Z(_12295_));
 MUX2_X1 _18209_ (.A(_00663_),
    .B(_00665_),
    .S(_12194_),
    .Z(_12296_));
 MUX2_X1 _18210_ (.A(_12295_),
    .B(_12296_),
    .S(_11955_),
    .Z(_12297_));
 MUX2_X1 _18211_ (.A(_12294_),
    .B(_12297_),
    .S(_12200_),
    .Z(_12298_));
 NOR2_X1 _18212_ (.A1(_12117_),
    .A2(_12298_),
    .ZN(_12299_));
 NOR3_X2 _18213_ (.A1(_11991_),
    .A2(_12291_),
    .A3(_12299_),
    .ZN(_12300_));
 MUX2_X1 _18214_ (.A(_00682_),
    .B(_00684_),
    .S(_12204_),
    .Z(_12301_));
 MUX2_X1 _18215_ (.A(_00683_),
    .B(_00685_),
    .S(_12204_),
    .Z(_12302_));
 MUX2_X1 _18216_ (.A(_12301_),
    .B(_12302_),
    .S(_12207_),
    .Z(_12303_));
 MUX2_X1 _18217_ (.A(_00674_),
    .B(_00676_),
    .S(_12204_),
    .Z(_12304_));
 MUX2_X1 _18218_ (.A(_00675_),
    .B(_00677_),
    .S(_12204_),
    .Z(_12305_));
 MUX2_X1 _18219_ (.A(_12304_),
    .B(_12305_),
    .S(_12207_),
    .Z(_12306_));
 MUX2_X1 _18220_ (.A(_12303_),
    .B(_12306_),
    .S(_12029_),
    .Z(_12307_));
 MUX2_X1 _18221_ (.A(_00686_),
    .B(_00688_),
    .S(_12204_),
    .Z(_12308_));
 MUX2_X1 _18222_ (.A(_00687_),
    .B(_00689_),
    .S(_12204_),
    .Z(_12309_));
 MUX2_X1 _18223_ (.A(_12308_),
    .B(_12309_),
    .S(_12207_),
    .Z(_12310_));
 MUX2_X1 _18224_ (.A(_00678_),
    .B(_00680_),
    .S(_12204_),
    .Z(_12311_));
 MUX2_X1 _18225_ (.A(_00679_),
    .B(_00681_),
    .S(_12021_),
    .Z(_12312_));
 MUX2_X1 _18226_ (.A(_12311_),
    .B(_12312_),
    .S(_12207_),
    .Z(_12313_));
 MUX2_X1 _18227_ (.A(_12310_),
    .B(_12313_),
    .S(_12029_),
    .Z(_12314_));
 MUX2_X1 _18228_ (.A(_12307_),
    .B(_12314_),
    .S(_11989_),
    .Z(_12315_));
 AOI21_X4 _18229_ (.A(_12300_),
    .B1(_11992_),
    .B2(_12315_),
    .ZN(_12316_));
 OAI221_X2 _18230_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12281_),
    .C1(_12316_),
    .C2(_11995_),
    .ZN(_15969_));
 INV_X1 _18231_ (.A(_15969_),
    .ZN(_15965_));
 BUF_X4 _18232_ (.A(_11639_),
    .Z(_12317_));
 MUX2_X1 _18233_ (.A(_00686_),
    .B(_00688_),
    .S(_12317_),
    .Z(_12318_));
 MUX2_X1 _18234_ (.A(_00687_),
    .B(_00689_),
    .S(_12317_),
    .Z(_12319_));
 MUX2_X1 _18235_ (.A(_12318_),
    .B(_12319_),
    .S(_10627_),
    .Z(_12320_));
 MUX2_X1 _18236_ (.A(_00678_),
    .B(_00680_),
    .S(_12317_),
    .Z(_12321_));
 MUX2_X1 _18237_ (.A(_00679_),
    .B(_00681_),
    .S(_12317_),
    .Z(_12322_));
 MUX2_X1 _18238_ (.A(_12321_),
    .B(_12322_),
    .S(_10627_),
    .Z(_12323_));
 MUX2_X1 _18239_ (.A(_12320_),
    .B(_12323_),
    .S(_10828_),
    .Z(_12324_));
 MUX2_X1 _18240_ (.A(_00682_),
    .B(_00684_),
    .S(_12317_),
    .Z(_12325_));
 MUX2_X1 _18241_ (.A(_00683_),
    .B(_00685_),
    .S(_12317_),
    .Z(_12326_));
 MUX2_X1 _18242_ (.A(_12325_),
    .B(_12326_),
    .S(_10627_),
    .Z(_12327_));
 MUX2_X1 _18243_ (.A(_00674_),
    .B(_00676_),
    .S(_12317_),
    .Z(_12328_));
 MUX2_X1 _18244_ (.A(_00675_),
    .B(_00677_),
    .S(_12317_),
    .Z(_12329_));
 MUX2_X1 _18245_ (.A(_12328_),
    .B(_12329_),
    .S(_10627_),
    .Z(_12330_));
 MUX2_X1 _18246_ (.A(_12327_),
    .B(_12330_),
    .S(_10828_),
    .Z(_12331_));
 MUX2_X1 _18247_ (.A(_12324_),
    .B(_12331_),
    .S(_10608_),
    .Z(_12332_));
 MUX2_X1 _18248_ (.A(_00670_),
    .B(_00672_),
    .S(_11597_),
    .Z(_12333_));
 MUX2_X1 _18249_ (.A(_00671_),
    .B(_00673_),
    .S(_11597_),
    .Z(_12334_));
 MUX2_X1 _18250_ (.A(_12333_),
    .B(_12334_),
    .S(_10797_),
    .Z(_12335_));
 NAND2_X1 _18251_ (.A1(_11533_),
    .A2(_12335_),
    .ZN(_12336_));
 MUX2_X1 _18252_ (.A(_00662_),
    .B(_00664_),
    .S(_11597_),
    .Z(_12337_));
 MUX2_X1 _18253_ (.A(_00663_),
    .B(_00665_),
    .S(_11597_),
    .Z(_12338_));
 MUX2_X1 _18254_ (.A(_12337_),
    .B(_12338_),
    .S(_10797_),
    .Z(_12339_));
 NAND2_X1 _18255_ (.A1(_10570_),
    .A2(_12339_),
    .ZN(_12340_));
 NAND3_X2 _18256_ (.A1(_10752_),
    .A2(_12336_),
    .A3(_12340_),
    .ZN(_12341_));
 NAND2_X1 _18257_ (.A1(_10602_),
    .A2(_00661_),
    .ZN(_12342_));
 OAI21_X1 _18258_ (.A(_12342_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .B2(_10589_),
    .ZN(_12343_));
 OAI221_X2 _18259_ (.A(_10570_),
    .B1(_00660_),
    .B2(_10757_),
    .C1(_12343_),
    .C2(_10581_),
    .ZN(_12344_));
 MUX2_X1 _18260_ (.A(_00666_),
    .B(_00668_),
    .S(_10600_),
    .Z(_12345_));
 MUX2_X1 _18261_ (.A(_00667_),
    .B(_00669_),
    .S(_10600_),
    .Z(_12346_));
 MUX2_X1 _18262_ (.A(_12345_),
    .B(_12346_),
    .S(_10628_),
    .Z(_12347_));
 AOI21_X1 _18263_ (.A(_11676_),
    .B1(_10766_),
    .B2(_12347_),
    .ZN(_12348_));
 AOI21_X2 _18264_ (.A(_10749_),
    .B1(_12344_),
    .B2(_12348_),
    .ZN(_12349_));
 AOI22_X4 _18265_ (.A1(_10750_),
    .A2(_12332_),
    .B1(_12341_),
    .B2(_12349_),
    .ZN(_12350_));
 NAND2_X1 _18266_ (.A1(_11596_),
    .A2(_12350_),
    .ZN(_12351_));
 INV_X1 _18267_ (.A(\cs_registers_i.pc_id_i[16] ),
    .ZN(_12352_));
 NOR2_X1 _18268_ (.A1(_12352_),
    .A2(_10668_),
    .ZN(_12353_));
 AOI22_X2 _18269_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(_10397_),
    .B1(_10683_),
    .B2(_12353_),
    .ZN(_12354_));
 NAND2_X2 _18270_ (.A1(_12351_),
    .A2(_12354_),
    .ZN(_15964_));
 INV_X4 _18271_ (.A(_15964_),
    .ZN(_15968_));
 NOR3_X1 _18272_ (.A1(_10610_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12355_));
 BUF_X32 _18273_ (.A(_11937_),
    .Z(_12356_));
 MUX2_X1 _18274_ (.A(_00713_),
    .B(_00715_),
    .S(_12356_),
    .Z(_12357_));
 MUX2_X1 _18275_ (.A(_00714_),
    .B(_00716_),
    .S(net402),
    .Z(_12358_));
 BUF_X4 _18276_ (.A(_11933_),
    .Z(_12359_));
 MUX2_X1 _18277_ (.A(_12357_),
    .B(_12358_),
    .S(_12359_),
    .Z(_12360_));
 MUX2_X1 _18278_ (.A(_00705_),
    .B(_00707_),
    .S(_12356_),
    .Z(_12361_));
 MUX2_X1 _18279_ (.A(_00706_),
    .B(_00708_),
    .S(_12356_),
    .Z(_12362_));
 MUX2_X1 _18280_ (.A(_12361_),
    .B(_12362_),
    .S(_12359_),
    .Z(_12363_));
 MUX2_X1 _18281_ (.A(_12360_),
    .B(_12363_),
    .S(_12005_),
    .Z(_12364_));
 NOR2_X4 _18282_ (.A1(_12364_),
    .A2(_11989_),
    .ZN(_12365_));
 MUX2_X1 _18283_ (.A(_00717_),
    .B(_00719_),
    .S(_11962_),
    .Z(_12366_));
 MUX2_X1 _18284_ (.A(_00718_),
    .B(_00720_),
    .S(_11962_),
    .Z(_12367_));
 MUX2_X1 _18285_ (.A(_12366_),
    .B(_12367_),
    .S(_11964_),
    .Z(_12368_));
 MUX2_X1 _18286_ (.A(_00709_),
    .B(_00711_),
    .S(_11962_),
    .Z(_12369_));
 MUX2_X1 _18287_ (.A(_00710_),
    .B(_00712_),
    .S(_11962_),
    .Z(_12370_));
 MUX2_X1 _18288_ (.A(_12369_),
    .B(_12370_),
    .S(_11964_),
    .Z(_12371_));
 MUX2_X1 _18289_ (.A(_12368_),
    .B(_12371_),
    .S(_11969_),
    .Z(_12372_));
 NOR2_X4 _18290_ (.A1(_11959_),
    .A2(_12372_),
    .ZN(_12373_));
 NOR3_X4 _18291_ (.A1(_12365_),
    .A2(_10474_),
    .A3(_12373_),
    .ZN(_12374_));
 MUX2_X1 _18292_ (.A(_00701_),
    .B(_00703_),
    .S(_12129_),
    .Z(_12375_));
 MUX2_X1 _18293_ (.A(_00702_),
    .B(_00704_),
    .S(_12129_),
    .Z(_12376_));
 MUX2_X1 _18294_ (.A(_12375_),
    .B(_12376_),
    .S(_12000_),
    .Z(_12377_));
 MUX2_X1 _18295_ (.A(_00693_),
    .B(_00695_),
    .S(_12129_),
    .Z(_12378_));
 MUX2_X1 _18296_ (.A(_00694_),
    .B(_00696_),
    .S(_12129_),
    .Z(_12379_));
 MUX2_X1 _18297_ (.A(_12378_),
    .B(_12379_),
    .S(_12207_),
    .Z(_12380_));
 MUX2_X1 _18298_ (.A(_12377_),
    .B(_12380_),
    .S(_12029_),
    .Z(_12381_));
 NOR2_X4 _18299_ (.A1(_12381_),
    .A2(_11959_),
    .ZN(_12382_));
 INV_X1 _18300_ (.A(_00691_),
    .ZN(_12383_));
 NOR2_X1 _18301_ (.A1(_11939_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .ZN(_12384_));
 AOI21_X1 _18302_ (.A(_12384_),
    .B1(_00692_),
    .B2(_12037_),
    .ZN(_12385_));
 AOI221_X1 _18303_ (.A(_11948_),
    .B1(_12383_),
    .B2(_11949_),
    .C1(_12385_),
    .C2(_11956_),
    .ZN(_12386_));
 MUX2_X1 _18304_ (.A(_00697_),
    .B(_00699_),
    .S(_12037_),
    .Z(_12387_));
 MUX2_X1 _18305_ (.A(_00698_),
    .B(_00700_),
    .S(_12037_),
    .Z(_12388_));
 MUX2_X1 _18306_ (.A(_12387_),
    .B(_12388_),
    .S(_11935_),
    .Z(_12389_));
 AOI21_X2 _18307_ (.A(_12386_),
    .B1(_12389_),
    .B2(_12041_),
    .ZN(_12390_));
 AOI21_X4 _18308_ (.A(_12382_),
    .B1(_12390_),
    .B2(_11959_),
    .ZN(_12391_));
 AOI21_X4 _18309_ (.A(_12374_),
    .B1(_10474_),
    .B2(_12391_),
    .ZN(_12392_));
 OAI221_X2 _18310_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12355_),
    .C1(_12392_),
    .C2(_11995_),
    .ZN(_15977_));
 INV_X1 _18311_ (.A(_15977_),
    .ZN(_15973_));
 MUX2_X1 _18312_ (.A(_00697_),
    .B(_00699_),
    .S(_11874_),
    .Z(_12393_));
 MUX2_X1 _18313_ (.A(_00698_),
    .B(_00700_),
    .S(_11874_),
    .Z(_12394_));
 MUX2_X1 _18314_ (.A(_12393_),
    .B(_12394_),
    .S(_11877_),
    .Z(_12395_));
 NOR2_X1 _18315_ (.A1(_10587_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .ZN(_12396_));
 AOI21_X1 _18316_ (.A(_12396_),
    .B1(_00692_),
    .B2(_11547_),
    .ZN(_12397_));
 AOI22_X1 _18317_ (.A1(_12383_),
    .A2(_10822_),
    .B1(_12397_),
    .B2(_10628_),
    .ZN(_12398_));
 MUX2_X1 _18318_ (.A(_12395_),
    .B(_12398_),
    .S(_11358_),
    .Z(_12399_));
 MUX2_X1 _18319_ (.A(_00709_),
    .B(_00711_),
    .S(_11363_),
    .Z(_12400_));
 MUX2_X1 _18320_ (.A(_00710_),
    .B(_00712_),
    .S(_11363_),
    .Z(_12401_));
 MUX2_X1 _18321_ (.A(_12400_),
    .B(_12401_),
    .S(_11366_),
    .Z(_12402_));
 NAND2_X1 _18322_ (.A1(_10778_),
    .A2(_12402_),
    .ZN(_12403_));
 MUX2_X1 _18323_ (.A(_00705_),
    .B(_00706_),
    .S(_11877_),
    .Z(_12404_));
 AOI21_X1 _18324_ (.A(_10575_),
    .B1(_10785_),
    .B2(_12404_),
    .ZN(_12405_));
 MUX2_X1 _18325_ (.A(_00707_),
    .B(_00708_),
    .S(_11877_),
    .Z(_12406_));
 NAND2_X1 _18326_ (.A1(_10794_),
    .A2(_12406_),
    .ZN(_12407_));
 NAND3_X1 _18327_ (.A1(_12403_),
    .A2(_12405_),
    .A3(_12407_),
    .ZN(_12408_));
 MUX2_X1 _18328_ (.A(_00713_),
    .B(_00714_),
    .S(_10627_),
    .Z(_12409_));
 NOR3_X1 _18329_ (.A1(_10589_),
    .A2(_10751_),
    .A3(_12409_),
    .ZN(_12410_));
 MUX2_X1 _18330_ (.A(_00715_),
    .B(_00716_),
    .S(_11375_),
    .Z(_12411_));
 NOR3_X1 _18331_ (.A1(_10632_),
    .A2(_10832_),
    .A3(_12411_),
    .ZN(_12412_));
 MUX2_X1 _18332_ (.A(_00717_),
    .B(_00718_),
    .S(_10861_),
    .Z(_12413_));
 MUX2_X1 _18333_ (.A(_00719_),
    .B(_00720_),
    .S(_10861_),
    .Z(_12414_));
 MUX2_X1 _18334_ (.A(_12413_),
    .B(_12414_),
    .S(_11597_),
    .Z(_12415_));
 OAI21_X1 _18335_ (.A(_10765_),
    .B1(_12415_),
    .B2(_11775_),
    .ZN(_12416_));
 NOR3_X1 _18336_ (.A1(_12410_),
    .A2(_12412_),
    .A3(_12416_),
    .ZN(_12417_));
 MUX2_X1 _18337_ (.A(_00701_),
    .B(_00703_),
    .S(_10619_),
    .Z(_12418_));
 MUX2_X1 _18338_ (.A(_00702_),
    .B(_00704_),
    .S(_10619_),
    .Z(_12419_));
 MUX2_X1 _18339_ (.A(_12418_),
    .B(_12419_),
    .S(_10796_),
    .Z(_12420_));
 MUX2_X1 _18340_ (.A(_00693_),
    .B(_00695_),
    .S(_11568_),
    .Z(_12421_));
 MUX2_X1 _18341_ (.A(_00694_),
    .B(_00696_),
    .S(_11568_),
    .Z(_12422_));
 MUX2_X1 _18342_ (.A(_12421_),
    .B(_12422_),
    .S(_10796_),
    .Z(_12423_));
 MUX2_X1 _18343_ (.A(_12420_),
    .B(_12423_),
    .S(_10828_),
    .Z(_12424_));
 OAI222_X2 _18344_ (.A1(_10831_),
    .A2(_12399_),
    .B1(_12408_),
    .B2(_12417_),
    .C1(_12424_),
    .C2(_10855_),
    .ZN(_12425_));
 NAND2_X1 _18345_ (.A1(_10816_),
    .A2(_12425_),
    .ZN(_12426_));
 AND2_X1 _18346_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_10563_),
    .ZN(_12427_));
 AOI22_X2 _18347_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(_11632_),
    .B1(_10870_),
    .B2(_12427_),
    .ZN(_12428_));
 NAND2_X2 _18348_ (.A1(_12426_),
    .A2(_12428_),
    .ZN(_15972_));
 INV_X2 _18349_ (.A(_15972_),
    .ZN(_15976_));
 BUF_X2 _18350_ (.A(_15438_),
    .Z(_12429_));
 INV_X1 _18351_ (.A(_15433_),
    .ZN(_12430_));
 INV_X1 _18352_ (.A(_12268_),
    .ZN(_12431_));
 AOI221_X2 _18353_ (.A(_15429_),
    .B1(_12261_),
    .B2(_12431_),
    .C1(_15425_),
    .C2(_15430_),
    .ZN(_12432_));
 BUF_X1 _18354_ (.A(_15434_),
    .Z(_12433_));
 INV_X1 _18355_ (.A(_12433_),
    .ZN(_12434_));
 OAI21_X2 _18356_ (.A(_12430_),
    .B1(_12432_),
    .B2(_12434_),
    .ZN(_12435_));
 NOR3_X2 _18357_ (.A1(_12434_),
    .A2(_12267_),
    .A3(_12268_),
    .ZN(_12436_));
 AOI21_X4 _18358_ (.A(_12435_),
    .B1(_11910_),
    .B2(_12436_),
    .ZN(_12437_));
 XNOR2_X2 _18359_ (.A(_12429_),
    .B(_12437_),
    .ZN(\alu_adder_result_ex[17] ));
 AOI21_X1 _18360_ (.A(_15429_),
    .B1(_15425_),
    .B2(_15430_),
    .ZN(_12438_));
 OAI21_X1 _18361_ (.A(_12081_),
    .B1(_12097_),
    .B2(_12096_),
    .ZN(_12439_));
 AOI21_X1 _18362_ (.A(_15421_),
    .B1(_12439_),
    .B2(_12079_),
    .ZN(_12440_));
 NAND2_X1 _18363_ (.A1(_12087_),
    .A2(_12269_),
    .ZN(_12441_));
 OAI221_X2 _18364_ (.A(_12438_),
    .B1(_12440_),
    .B2(_12268_),
    .C1(_12441_),
    .C2(_11850_),
    .ZN(_12442_));
 NAND3_X1 _18365_ (.A1(_11839_),
    .A2(_12087_),
    .A3(_12269_),
    .ZN(_12443_));
 AOI211_X2 _18366_ (.A(_11854_),
    .B(_12443_),
    .C1(_11858_),
    .C2(_11918_),
    .ZN(_12444_));
 OAI21_X1 _18367_ (.A(_12433_),
    .B1(_12442_),
    .B2(_12444_),
    .ZN(_12445_));
 OR3_X1 _18368_ (.A1(_12433_),
    .A2(_12442_),
    .A3(_12444_),
    .ZN(_12446_));
 AND2_X1 _18369_ (.A1(_12445_),
    .A2(_12446_),
    .ZN(_12447_));
 BUF_X4 _18370_ (.A(_12447_),
    .Z(\alu_adder_result_ex[16] ));
 NOR3_X1 _18371_ (.A1(_10571_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12448_));
 CLKBUF_X3 _18372_ (.A(_10436_),
    .Z(_12449_));
 MUX2_X1 _18373_ (.A(_00728_),
    .B(_00730_),
    .S(_11952_),
    .Z(_12450_));
 MUX2_X1 _18374_ (.A(_00729_),
    .B(_00731_),
    .S(_11952_),
    .Z(_12451_));
 MUX2_X1 _18375_ (.A(_12450_),
    .B(_12451_),
    .S(_11975_),
    .Z(_12452_));
 NAND2_X1 _18376_ (.A1(_12041_),
    .A2(_12452_),
    .ZN(_12453_));
 NAND2_X1 _18377_ (.A1(_12037_),
    .A2(_00723_),
    .ZN(_12454_));
 OAI21_X1 _18378_ (.A(_12454_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B2(_12034_),
    .ZN(_12455_));
 OAI221_X1 _18379_ (.A(_12005_),
    .B1(_00722_),
    .B2(_10716_),
    .C1(_12455_),
    .C2(_11942_),
    .ZN(_12456_));
 AND3_X1 _18380_ (.A1(_12449_),
    .A2(_12453_),
    .A3(_12456_),
    .ZN(_12457_));
 MUX2_X1 _18381_ (.A(_00732_),
    .B(_00734_),
    .S(_12194_),
    .Z(_12458_));
 MUX2_X1 _18382_ (.A(_00733_),
    .B(_00735_),
    .S(_11960_),
    .Z(_12459_));
 MUX2_X1 _18383_ (.A(_12458_),
    .B(_12459_),
    .S(_11964_),
    .Z(_12460_));
 MUX2_X1 _18384_ (.A(_00724_),
    .B(_00726_),
    .S(_11960_),
    .Z(_12461_));
 MUX2_X1 _18385_ (.A(_00725_),
    .B(_00727_),
    .S(_11960_),
    .Z(_12462_));
 MUX2_X1 _18386_ (.A(_12461_),
    .B(_12462_),
    .S(_11964_),
    .Z(_12463_));
 MUX2_X1 _18387_ (.A(_12460_),
    .B(_12463_),
    .S(_12200_),
    .Z(_12464_));
 NOR2_X1 _18388_ (.A1(_12117_),
    .A2(_12464_),
    .ZN(_12465_));
 NOR3_X2 _18389_ (.A1(_11991_),
    .A2(_12457_),
    .A3(_12465_),
    .ZN(_12466_));
 MUX2_X1 _18390_ (.A(_00744_),
    .B(_00746_),
    .S(_12023_),
    .Z(_12467_));
 MUX2_X1 _18391_ (.A(_00745_),
    .B(_00747_),
    .S(_12023_),
    .Z(_12468_));
 MUX2_X1 _18392_ (.A(_12467_),
    .B(_12468_),
    .S(_11934_),
    .Z(_12469_));
 MUX2_X1 _18393_ (.A(_00736_),
    .B(_00738_),
    .S(_12023_),
    .Z(_12470_));
 MUX2_X1 _18394_ (.A(_00737_),
    .B(_00739_),
    .S(_12023_),
    .Z(_12471_));
 MUX2_X1 _18395_ (.A(_12470_),
    .B(_12471_),
    .S(_11934_),
    .Z(_12472_));
 MUX2_X1 _18396_ (.A(_12469_),
    .B(_12472_),
    .S(_12029_),
    .Z(_12473_));
 MUX2_X1 _18397_ (.A(_00748_),
    .B(_00750_),
    .S(_12023_),
    .Z(_12474_));
 MUX2_X1 _18398_ (.A(_00749_),
    .B(_00751_),
    .S(_11952_),
    .Z(_12475_));
 MUX2_X1 _18399_ (.A(_12474_),
    .B(_12475_),
    .S(_11975_),
    .Z(_12476_));
 MUX2_X1 _18400_ (.A(_00740_),
    .B(_00742_),
    .S(_12023_),
    .Z(_12477_));
 MUX2_X1 _18401_ (.A(_00741_),
    .B(_00743_),
    .S(_11952_),
    .Z(_12478_));
 MUX2_X1 _18402_ (.A(_12477_),
    .B(_12478_),
    .S(_11975_),
    .Z(_12479_));
 MUX2_X1 _18403_ (.A(_12476_),
    .B(_12479_),
    .S(_12029_),
    .Z(_12480_));
 MUX2_X1 _18404_ (.A(_12473_),
    .B(_12480_),
    .S(_11989_),
    .Z(_12481_));
 AOI21_X4 _18405_ (.A(_12466_),
    .B1(_12481_),
    .B2(_11992_),
    .ZN(_12482_));
 OAI221_X2 _18406_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12448_),
    .C1(_12482_),
    .C2(_11995_),
    .ZN(_15980_));
 INV_X1 _18407_ (.A(_15980_),
    .ZN(_15984_));
 NAND2_X1 _18408_ (.A1(_10602_),
    .A2(_00723_),
    .ZN(_12483_));
 OAI21_X1 _18409_ (.A(_12483_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B2(_10622_),
    .ZN(_12484_));
 OAI221_X1 _18410_ (.A(_10783_),
    .B1(_00722_),
    .B2(_10757_),
    .C1(_12484_),
    .C2(_10581_),
    .ZN(_12485_));
 MUX2_X1 _18411_ (.A(_00736_),
    .B(_00738_),
    .S(_10620_),
    .Z(_12486_));
 MUX2_X1 _18412_ (.A(_00737_),
    .B(_00739_),
    .S(_10620_),
    .Z(_12487_));
 MUX2_X1 _18413_ (.A(_12486_),
    .B(_12487_),
    .S(_10788_),
    .Z(_12488_));
 AOI21_X1 _18414_ (.A(_11437_),
    .B1(_12488_),
    .B2(_10749_),
    .ZN(_12489_));
 NAND2_X1 _18415_ (.A1(_12485_),
    .A2(_12489_),
    .ZN(_12490_));
 MUX2_X1 _18416_ (.A(_00744_),
    .B(_00746_),
    .S(_11874_),
    .Z(_12491_));
 MUX2_X1 _18417_ (.A(_00745_),
    .B(_00747_),
    .S(_11874_),
    .Z(_12492_));
 MUX2_X1 _18418_ (.A(_12491_),
    .B(_12492_),
    .S(_11877_),
    .Z(_12493_));
 MUX2_X1 _18419_ (.A(_00728_),
    .B(_00730_),
    .S(_11874_),
    .Z(_12494_));
 MUX2_X1 _18420_ (.A(_00729_),
    .B(_00731_),
    .S(_11874_),
    .Z(_12495_));
 MUX2_X1 _18421_ (.A(_12494_),
    .B(_12495_),
    .S(_11877_),
    .Z(_12496_));
 MUX2_X1 _18422_ (.A(_12493_),
    .B(_12496_),
    .S(_10575_),
    .Z(_12497_));
 BUF_X4 _18423_ (.A(_11655_),
    .Z(_12498_));
 MUX2_X1 _18424_ (.A(_00748_),
    .B(_00750_),
    .S(_12498_),
    .Z(_12499_));
 MUX2_X1 _18425_ (.A(_00749_),
    .B(_00751_),
    .S(_12498_),
    .Z(_12500_));
 MUX2_X1 _18426_ (.A(_12499_),
    .B(_12500_),
    .S(_10843_),
    .Z(_12501_));
 MUX2_X1 _18427_ (.A(_00732_),
    .B(_00734_),
    .S(_12498_),
    .Z(_12502_));
 MUX2_X1 _18428_ (.A(_00733_),
    .B(_00735_),
    .S(_12498_),
    .Z(_12503_));
 MUX2_X1 _18429_ (.A(_12502_),
    .B(_12503_),
    .S(_10843_),
    .Z(_12504_));
 MUX2_X1 _18430_ (.A(_12501_),
    .B(_12504_),
    .S(_10574_),
    .Z(_12505_));
 MUX2_X1 _18431_ (.A(_00740_),
    .B(_00742_),
    .S(_12498_),
    .Z(_12506_));
 MUX2_X1 _18432_ (.A(_00741_),
    .B(_00743_),
    .S(_12498_),
    .Z(_12507_));
 MUX2_X1 _18433_ (.A(_12506_),
    .B(_12507_),
    .S(_10839_),
    .Z(_12508_));
 MUX2_X1 _18434_ (.A(_00724_),
    .B(_00726_),
    .S(_12498_),
    .Z(_12509_));
 MUX2_X1 _18435_ (.A(_00725_),
    .B(_00727_),
    .S(_10791_),
    .Z(_12510_));
 MUX2_X1 _18436_ (.A(_12509_),
    .B(_12510_),
    .S(_10839_),
    .Z(_12511_));
 MUX2_X1 _18437_ (.A(_12508_),
    .B(_12511_),
    .S(_10574_),
    .Z(_12512_));
 MUX2_X1 _18438_ (.A(_12505_),
    .B(_12512_),
    .S(_11358_),
    .Z(_12513_));
 OAI221_X2 _18439_ (.A(_12490_),
    .B1(_12497_),
    .B2(_11453_),
    .C1(_12513_),
    .C2(_10609_),
    .ZN(_12514_));
 NAND2_X1 _18440_ (.A1(_11596_),
    .A2(_12514_),
    .ZN(_12515_));
 AND2_X1 _18441_ (.A1(\cs_registers_i.pc_id_i[18] ),
    .A2(_11593_),
    .ZN(_12516_));
 AOI22_X4 _18442_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(_10741_),
    .B1(_10870_),
    .B2(_12516_),
    .ZN(_12517_));
 NAND2_X4 _18443_ (.A1(_12515_),
    .A2(_12517_),
    .ZN(_15985_));
 INV_X2 _18444_ (.A(_15985_),
    .ZN(_15981_));
 NOR3_X1 _18445_ (.A1(_10576_),
    .A2(_10398_),
    .A3(_11926_),
    .ZN(_12518_));
 MUX2_X1 _18446_ (.A(_00775_),
    .B(_00777_),
    .S(_11997_),
    .Z(_12519_));
 MUX2_X1 _18447_ (.A(_00776_),
    .B(_00778_),
    .S(_11997_),
    .Z(_12520_));
 MUX2_X1 _18448_ (.A(_12519_),
    .B(_12520_),
    .S(_12000_),
    .Z(_12521_));
 MUX2_X1 _18449_ (.A(_00767_),
    .B(_00769_),
    .S(_11997_),
    .Z(_12522_));
 MUX2_X1 _18450_ (.A(_00768_),
    .B(_00770_),
    .S(_11997_),
    .Z(_12523_));
 MUX2_X1 _18451_ (.A(_12522_),
    .B(_12523_),
    .S(_12000_),
    .Z(_12524_));
 MUX2_X1 _18452_ (.A(_12521_),
    .B(_12524_),
    .S(_12005_),
    .Z(_12525_));
 NOR2_X2 _18453_ (.A1(_11989_),
    .A2(_12525_),
    .ZN(_12526_));
 MUX2_X1 _18454_ (.A(_00779_),
    .B(_00781_),
    .S(_12008_),
    .Z(_12527_));
 MUX2_X1 _18455_ (.A(_00780_),
    .B(_00782_),
    .S(_12008_),
    .Z(_12528_));
 MUX2_X1 _18456_ (.A(_12527_),
    .B(_12528_),
    .S(_12012_),
    .Z(_12529_));
 MUX2_X1 _18457_ (.A(_00771_),
    .B(_00773_),
    .S(_12008_),
    .Z(_12530_));
 MUX2_X1 _18458_ (.A(_00772_),
    .B(_00774_),
    .S(_12010_),
    .Z(_12531_));
 MUX2_X1 _18459_ (.A(_12530_),
    .B(_12531_),
    .S(_12012_),
    .Z(_12532_));
 MUX2_X1 _18460_ (.A(_12529_),
    .B(_12532_),
    .S(_12017_),
    .Z(_12533_));
 NOR2_X4 _18461_ (.A1(_12533_),
    .A2(_11959_),
    .ZN(_12534_));
 NOR3_X4 _18462_ (.A1(_12534_),
    .A2(_12526_),
    .A3(_10474_),
    .ZN(_12535_));
 MUX2_X1 _18463_ (.A(_00763_),
    .B(_00765_),
    .S(_12021_),
    .Z(_12536_));
 MUX2_X1 _18464_ (.A(_00764_),
    .B(_00766_),
    .S(_12021_),
    .Z(_12537_));
 MUX2_X1 _18465_ (.A(_12536_),
    .B(_12537_),
    .S(_11934_),
    .Z(_12538_));
 MUX2_X1 _18466_ (.A(_00755_),
    .B(_00757_),
    .S(_12021_),
    .Z(_12539_));
 MUX2_X1 _18467_ (.A(_00756_),
    .B(_00758_),
    .S(_12023_),
    .Z(_12540_));
 MUX2_X1 _18468_ (.A(_12539_),
    .B(_12540_),
    .S(_11934_),
    .Z(_12541_));
 MUX2_X1 _18469_ (.A(_12538_),
    .B(_12541_),
    .S(_12029_),
    .Z(_12542_));
 NOR2_X1 _18470_ (.A1(_11959_),
    .A2(_12542_),
    .ZN(_12543_));
 INV_X1 _18471_ (.A(_00753_),
    .ZN(_12544_));
 NOR2_X1 _18472_ (.A1(_11939_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .ZN(_12545_));
 AOI21_X1 _18473_ (.A(_12545_),
    .B1(_00754_),
    .B2(_12034_),
    .ZN(_12546_));
 AOI221_X1 _18474_ (.A(_11948_),
    .B1(_12544_),
    .B2(_11949_),
    .C1(_12546_),
    .C2(_11956_),
    .ZN(_12547_));
 MUX2_X1 _18475_ (.A(_00759_),
    .B(_00761_),
    .S(_12037_),
    .Z(_12548_));
 MUX2_X1 _18476_ (.A(_00760_),
    .B(_00762_),
    .S(_12037_),
    .Z(_12549_));
 MUX2_X1 _18477_ (.A(_12548_),
    .B(_12549_),
    .S(_11935_),
    .Z(_12550_));
 AOI21_X1 _18478_ (.A(_12547_),
    .B1(_12550_),
    .B2(_12041_),
    .ZN(_12551_));
 AOI21_X2 _18479_ (.A(_12543_),
    .B1(_12551_),
    .B2(_11959_),
    .ZN(_12552_));
 AOI21_X4 _18480_ (.A(_12535_),
    .B1(_12552_),
    .B2(_10474_),
    .ZN(_12553_));
 OAI221_X2 _18481_ (.A(_11922_),
    .B1(_11925_),
    .B2(_12518_),
    .C1(_12553_),
    .C2(_11995_),
    .ZN(_15993_));
 INV_X1 _18482_ (.A(_15993_),
    .ZN(_15989_));
 MUX2_X1 _18483_ (.A(_00767_),
    .B(_00768_),
    .S(_10593_),
    .Z(_12554_));
 AOI21_X1 _18484_ (.A(_10573_),
    .B1(_10785_),
    .B2(_12554_),
    .ZN(_12555_));
 MUX2_X1 _18485_ (.A(_00769_),
    .B(_00770_),
    .S(_10593_),
    .Z(_12556_));
 NAND3_X1 _18486_ (.A1(_10614_),
    .A2(_10792_),
    .A3(_12556_),
    .ZN(_12557_));
 NAND2_X1 _18487_ (.A1(_12555_),
    .A2(_12557_),
    .ZN(_12558_));
 MUX2_X1 _18488_ (.A(_00771_),
    .B(_00773_),
    .S(_11545_),
    .Z(_12559_));
 MUX2_X1 _18489_ (.A(_00772_),
    .B(_00774_),
    .S(_11545_),
    .Z(_12560_));
 MUX2_X1 _18490_ (.A(_12559_),
    .B(_12560_),
    .S(_10594_),
    .Z(_12561_));
 MUX2_X1 _18491_ (.A(_00777_),
    .B(_00778_),
    .S(_10577_),
    .Z(_12562_));
 MUX2_X1 _18492_ (.A(_00775_),
    .B(_00776_),
    .S(_10577_),
    .Z(_12563_));
 MUX2_X1 _18493_ (.A(_12562_),
    .B(_12563_),
    .S(_10632_),
    .Z(_12564_));
 MUX2_X1 _18494_ (.A(_00781_),
    .B(_00782_),
    .S(_10577_),
    .Z(_12565_));
 MUX2_X1 _18495_ (.A(_00779_),
    .B(_00780_),
    .S(_10577_),
    .Z(_12566_));
 MUX2_X1 _18496_ (.A(_12565_),
    .B(_12566_),
    .S(_10632_),
    .Z(_12567_));
 MUX2_X1 _18497_ (.A(_12564_),
    .B(_12567_),
    .S(_10606_),
    .Z(_12568_));
 AOI221_X2 _18498_ (.A(_12558_),
    .B1(_12561_),
    .B2(_10778_),
    .C1(_10766_),
    .C2(_12568_),
    .ZN(_12569_));
 MUX2_X1 _18499_ (.A(_00759_),
    .B(_00761_),
    .S(_11546_),
    .Z(_12570_));
 NOR2_X1 _18500_ (.A1(_10628_),
    .A2(_12570_),
    .ZN(_12571_));
 MUX2_X1 _18501_ (.A(_00760_),
    .B(_00762_),
    .S(_11454_),
    .Z(_12572_));
 NOR2_X1 _18502_ (.A1(_10580_),
    .A2(_12572_),
    .ZN(_12573_));
 NOR3_X1 _18503_ (.A1(_11358_),
    .A2(_12571_),
    .A3(_12573_),
    .ZN(_12574_));
 NOR2_X1 _18504_ (.A1(_11874_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .ZN(_12575_));
 AOI21_X1 _18505_ (.A(_12575_),
    .B1(_00754_),
    .B2(_10587_),
    .ZN(_12576_));
 AOI221_X1 _18506_ (.A(_10765_),
    .B1(_12544_),
    .B2(_10822_),
    .C1(_12576_),
    .C2(_11877_),
    .ZN(_12577_));
 MUX2_X1 _18507_ (.A(_00763_),
    .B(_00765_),
    .S(_11874_),
    .Z(_12578_));
 NOR2_X1 _18508_ (.A1(_11535_),
    .A2(_12578_),
    .ZN(_12579_));
 MUX2_X1 _18509_ (.A(_00764_),
    .B(_00766_),
    .S(_11874_),
    .Z(_12580_));
 NOR2_X1 _18510_ (.A1(_10580_),
    .A2(_12580_),
    .ZN(_12581_));
 NOR3_X1 _18511_ (.A1(_10828_),
    .A2(_12579_),
    .A3(_12581_),
    .ZN(_12582_));
 MUX2_X1 _18512_ (.A(_00755_),
    .B(_00757_),
    .S(_11568_),
    .Z(_12583_));
 NOR2_X1 _18513_ (.A1(_10595_),
    .A2(_12583_),
    .ZN(_12584_));
 MUX2_X1 _18514_ (.A(_00756_),
    .B(_00758_),
    .S(_11568_),
    .Z(_12585_));
 NOR2_X1 _18515_ (.A1(_10580_),
    .A2(_12585_),
    .ZN(_12586_));
 NOR3_X1 _18516_ (.A1(_10765_),
    .A2(_12584_),
    .A3(_12586_),
    .ZN(_12587_));
 OAI33_X1 _18517_ (.A1(_10831_),
    .A2(_12574_),
    .A3(_12577_),
    .B1(_12582_),
    .B2(_12587_),
    .B3(_10855_),
    .ZN(_12588_));
 OR2_X4 _18518_ (.A1(_12569_),
    .A2(_12588_),
    .ZN(_12589_));
 BUF_X2 _18519_ (.A(\cs_registers_i.pc_id_i[19] ),
    .Z(_12590_));
 AND2_X1 _18520_ (.A1(_12590_),
    .A2(_11593_),
    .ZN(_12591_));
 AOI222_X2 _18521_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(_10741_),
    .B1(_10816_),
    .B2(_12589_),
    .C1(_12591_),
    .C2(_10870_),
    .ZN(_15992_));
 CLKBUF_X3 _18522_ (.A(_15446_),
    .Z(_12592_));
 BUF_X2 _18523_ (.A(_15442_),
    .Z(_12593_));
 INV_X1 _18524_ (.A(_12593_),
    .ZN(_12594_));
 INV_X1 _18525_ (.A(_15437_),
    .ZN(_12595_));
 OAI21_X1 _18526_ (.A(_12429_),
    .B1(_15433_),
    .B2(_12433_),
    .ZN(_12596_));
 AOI21_X2 _18527_ (.A(_12594_),
    .B1(_12595_),
    .B2(_12596_),
    .ZN(_12597_));
 AOI21_X2 _18528_ (.A(_15441_),
    .B1(_15437_),
    .B2(_12593_),
    .ZN(_12598_));
 NAND3_X2 _18529_ (.A1(_12430_),
    .A2(net448),
    .A3(_12598_),
    .ZN(_12599_));
 OAI22_X4 _18530_ (.A1(_15441_),
    .A2(_12597_),
    .B1(_12599_),
    .B2(_12270_),
    .ZN(_12600_));
 XNOR2_X2 _18531_ (.A(_12600_),
    .B(_12592_),
    .ZN(\alu_adder_result_ex[19] ));
 AND3_X1 _18532_ (.A1(_12433_),
    .A2(_12429_),
    .A3(_12269_),
    .ZN(_12601_));
 AND3_X1 _18533_ (.A1(_11902_),
    .A2(_11900_),
    .A3(_12601_),
    .ZN(_12602_));
 NAND2_X4 _18534_ (.A1(_11916_),
    .A2(_12602_),
    .ZN(_12603_));
 AND3_X2 _18535_ (.A1(_11839_),
    .A2(_12087_),
    .A3(_12601_),
    .ZN(_12604_));
 OAI211_X4 _18536_ (.A(_11501_),
    .B(_12604_),
    .C1(_11513_),
    .C2(_11862_),
    .ZN(_12605_));
 NAND3_X1 _18537_ (.A1(_11900_),
    .A2(_11901_),
    .A3(_12269_),
    .ZN(_12606_));
 AOI21_X1 _18538_ (.A(_12434_),
    .B1(_12432_),
    .B2(_12606_),
    .ZN(_12607_));
 OAI21_X2 _18539_ (.A(_12429_),
    .B1(_15433_),
    .B2(_12607_),
    .ZN(_12608_));
 AND2_X2 _18540_ (.A1(_12595_),
    .A2(_12608_),
    .ZN(_12609_));
 AND3_X4 _18541_ (.A1(_12603_),
    .A2(_12605_),
    .A3(_12609_),
    .ZN(_12610_));
 XNOR2_X2 _18542_ (.A(_12593_),
    .B(_12610_),
    .ZN(\alu_adder_result_ex[18] ));
 AOI21_X2 _18543_ (.A(_11923_),
    .B1(_11320_),
    .B2(_10928_),
    .ZN(_12611_));
 OAI21_X2 _18544_ (.A(_10317_),
    .B1(_12611_),
    .B2(_10398_),
    .ZN(_12612_));
 BUF_X2 _18545_ (.A(_12612_),
    .Z(_12613_));
 CLKBUF_X3 _18546_ (.A(_11162_),
    .Z(_12614_));
 AOI21_X1 _18547_ (.A(_12613_),
    .B1(_12614_),
    .B2(_11935_),
    .ZN(_12615_));
 MUX2_X1 _18548_ (.A(_00790_),
    .B(_00792_),
    .S(_11960_),
    .Z(_12616_));
 MUX2_X1 _18549_ (.A(_00791_),
    .B(_00793_),
    .S(_11960_),
    .Z(_12617_));
 MUX2_X1 _18550_ (.A(_12616_),
    .B(_12617_),
    .S(_11964_),
    .Z(_12618_));
 NAND2_X1 _18551_ (.A1(_11948_),
    .A2(_12618_),
    .ZN(_12619_));
 NAND2_X1 _18552_ (.A1(_11953_),
    .A2(_00785_),
    .ZN(_12620_));
 OAI21_X1 _18553_ (.A(_12620_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B2(_12037_),
    .ZN(_12621_));
 OAI221_X1 _18554_ (.A(_12124_),
    .B1(_00784_),
    .B2(_10716_),
    .C1(_12621_),
    .C2(_10697_),
    .ZN(_12622_));
 AND3_X1 _18555_ (.A1(_10436_),
    .A2(_12619_),
    .A3(_12622_),
    .ZN(_12623_));
 MUX2_X1 _18556_ (.A(_00794_),
    .B(_00796_),
    .S(_11951_),
    .Z(_12624_));
 MUX2_X1 _18557_ (.A(_00795_),
    .B(_00797_),
    .S(_11951_),
    .Z(_12625_));
 MUX2_X1 _18558_ (.A(_12624_),
    .B(_12625_),
    .S(_11933_),
    .Z(_12626_));
 MUX2_X1 _18559_ (.A(_00786_),
    .B(_00788_),
    .S(_11951_),
    .Z(_12627_));
 BUF_X4 _18560_ (.A(net357),
    .Z(_12628_));
 MUX2_X1 _18561_ (.A(_00787_),
    .B(_00789_),
    .S(_12628_),
    .Z(_12629_));
 BUF_X4 _18562_ (.A(_10466_),
    .Z(_12630_));
 MUX2_X1 _18563_ (.A(_12627_),
    .B(_12629_),
    .S(_12630_),
    .Z(_12631_));
 MUX2_X1 _18564_ (.A(_12626_),
    .B(_12631_),
    .S(_11931_),
    .Z(_12632_));
 NOR2_X1 _18565_ (.A1(_12449_),
    .A2(_12632_),
    .ZN(_12633_));
 NOR3_X2 _18566_ (.A1(_11928_),
    .A2(_12623_),
    .A3(_12633_),
    .ZN(_12634_));
 MUX2_X1 _18567_ (.A(_00806_),
    .B(_00808_),
    .S(_12194_),
    .Z(_12635_));
 MUX2_X1 _18568_ (.A(_00807_),
    .B(_00809_),
    .S(_12194_),
    .Z(_12636_));
 MUX2_X1 _18569_ (.A(_12635_),
    .B(_12636_),
    .S(_11955_),
    .Z(_12637_));
 MUX2_X1 _18570_ (.A(_00798_),
    .B(_00800_),
    .S(_12194_),
    .Z(_12638_));
 MUX2_X1 _18571_ (.A(_00799_),
    .B(_00801_),
    .S(_11960_),
    .Z(_12639_));
 MUX2_X1 _18572_ (.A(_12638_),
    .B(_12639_),
    .S(_11955_),
    .Z(_12640_));
 MUX2_X1 _18573_ (.A(_12637_),
    .B(_12640_),
    .S(_12200_),
    .Z(_12641_));
 MUX2_X1 _18574_ (.A(_00810_),
    .B(_00812_),
    .S(_12194_),
    .Z(_12642_));
 MUX2_X1 _18575_ (.A(_00811_),
    .B(_00813_),
    .S(_11960_),
    .Z(_12643_));
 MUX2_X1 _18576_ (.A(_12642_),
    .B(_12643_),
    .S(_11964_),
    .Z(_12644_));
 MUX2_X1 _18577_ (.A(_00802_),
    .B(_00804_),
    .S(_11960_),
    .Z(_12645_));
 MUX2_X1 _18578_ (.A(_00803_),
    .B(_00805_),
    .S(_11960_),
    .Z(_12646_));
 MUX2_X1 _18579_ (.A(_12645_),
    .B(_12646_),
    .S(_11964_),
    .Z(_12647_));
 MUX2_X1 _18580_ (.A(_12644_),
    .B(_12647_),
    .S(_12200_),
    .Z(_12648_));
 BUF_X4 _18581_ (.A(_10432_),
    .Z(_12649_));
 MUX2_X1 _18582_ (.A(_12641_),
    .B(_12648_),
    .S(_12649_),
    .Z(_12650_));
 AOI21_X4 _18583_ (.A(_12634_),
    .B1(_12650_),
    .B2(_11929_),
    .ZN(_12651_));
 OAI21_X1 _18584_ (.A(_11922_),
    .B1(_11995_),
    .B2(_12651_),
    .ZN(_12652_));
 NOR2_X2 _18585_ (.A1(_12615_),
    .A2(_12652_),
    .ZN(_16000_));
 MUX2_X1 _18586_ (.A(_00790_),
    .B(_00792_),
    .S(_11597_),
    .Z(_12653_));
 MUX2_X1 _18587_ (.A(_00791_),
    .B(_00793_),
    .S(_10614_),
    .Z(_12654_));
 MUX2_X1 _18588_ (.A(_12653_),
    .B(_12654_),
    .S(_10797_),
    .Z(_12655_));
 AOI21_X1 _18589_ (.A(_10831_),
    .B1(_12655_),
    .B2(_11533_),
    .ZN(_12656_));
 NAND2_X1 _18590_ (.A1(_10589_),
    .A2(_00785_),
    .ZN(_12657_));
 OAI21_X1 _18591_ (.A(_12657_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B2(_10622_),
    .ZN(_12658_));
 OAI22_X1 _18592_ (.A1(_00784_),
    .A2(_10758_),
    .B1(_12658_),
    .B2(_10581_),
    .ZN(_12659_));
 OAI21_X1 _18593_ (.A(_12656_),
    .B1(_12659_),
    .B2(_10767_),
    .ZN(_12660_));
 MUX2_X1 _18594_ (.A(_00806_),
    .B(_00808_),
    .S(_10823_),
    .Z(_12661_));
 MUX2_X1 _18595_ (.A(_00807_),
    .B(_00809_),
    .S(_10823_),
    .Z(_12662_));
 MUX2_X1 _18596_ (.A(_12661_),
    .B(_12662_),
    .S(_11535_),
    .Z(_12663_));
 MUX2_X1 _18597_ (.A(_00798_),
    .B(_00800_),
    .S(_10823_),
    .Z(_12664_));
 MUX2_X1 _18598_ (.A(_00799_),
    .B(_00801_),
    .S(_10823_),
    .Z(_12665_));
 MUX2_X1 _18599_ (.A(_12664_),
    .B(_12665_),
    .S(_11535_),
    .Z(_12666_));
 MUX2_X1 _18600_ (.A(_12663_),
    .B(_12666_),
    .S(_11358_),
    .Z(_12667_));
 MUX2_X1 _18601_ (.A(_00810_),
    .B(_00812_),
    .S(_11545_),
    .Z(_12668_));
 MUX2_X1 _18602_ (.A(_00811_),
    .B(_00813_),
    .S(_11614_),
    .Z(_12669_));
 MUX2_X1 _18603_ (.A(_12668_),
    .B(_12669_),
    .S(_10594_),
    .Z(_12670_));
 MUX2_X1 _18604_ (.A(_00802_),
    .B(_00804_),
    .S(_11614_),
    .Z(_12671_));
 MUX2_X1 _18605_ (.A(_00803_),
    .B(_00805_),
    .S(_11614_),
    .Z(_12672_));
 MUX2_X1 _18606_ (.A(_12671_),
    .B(_12672_),
    .S(_11375_),
    .Z(_12673_));
 MUX2_X1 _18607_ (.A(_12670_),
    .B(_12673_),
    .S(_10569_),
    .Z(_12674_));
 MUX2_X1 _18608_ (.A(_00794_),
    .B(_00796_),
    .S(_11614_),
    .Z(_12675_));
 MUX2_X1 _18609_ (.A(_00795_),
    .B(_00797_),
    .S(_11372_),
    .Z(_12676_));
 MUX2_X1 _18610_ (.A(_12675_),
    .B(_12676_),
    .S(_11375_),
    .Z(_12677_));
 MUX2_X1 _18611_ (.A(_00786_),
    .B(_00788_),
    .S(_11372_),
    .Z(_12678_));
 MUX2_X1 _18612_ (.A(_00787_),
    .B(_00789_),
    .S(_11372_),
    .Z(_12679_));
 MUX2_X1 _18613_ (.A(_12678_),
    .B(_12679_),
    .S(_11375_),
    .Z(_12680_));
 MUX2_X1 _18614_ (.A(_12677_),
    .B(_12680_),
    .S(_10569_),
    .Z(_12681_));
 MUX2_X1 _18615_ (.A(_12674_),
    .B(_12681_),
    .S(_10783_),
    .Z(_12682_));
 OAI221_X2 _18616_ (.A(_12660_),
    .B1(_12667_),
    .B2(_11371_),
    .C1(_10610_),
    .C2(_12682_),
    .ZN(_12683_));
 NAND2_X1 _18617_ (.A1(_11596_),
    .A2(net360),
    .ZN(_12684_));
 BUF_X2 _18618_ (.A(\cs_registers_i.pc_id_i[20] ),
    .Z(_12685_));
 AND2_X1 _18619_ (.A1(_12685_),
    .A2(_11593_),
    .ZN(_12686_));
 AOI22_X4 _18620_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(_10741_),
    .B1(_10683_),
    .B2(_12686_),
    .ZN(_12687_));
 NAND2_X4 _18621_ (.A1(_12684_),
    .A2(_12687_),
    .ZN(_16001_));
 INV_X2 _18622_ (.A(_16001_),
    .ZN(_15997_));
 AOI21_X1 _18623_ (.A(_12613_),
    .B1(_12614_),
    .B2(_12034_),
    .ZN(_12688_));
 BUF_X32 _18624_ (.A(net430),
    .Z(_12689_));
 MUX2_X1 _18625_ (.A(_00821_),
    .B(_00823_),
    .S(_12689_),
    .Z(_12690_));
 BUF_X32 _18626_ (.A(net326),
    .Z(_12691_));
 MUX2_X1 _18627_ (.A(_00822_),
    .B(_00824_),
    .S(_12691_),
    .Z(_12692_));
 BUF_X4 _18628_ (.A(_10466_),
    .Z(_12693_));
 MUX2_X1 _18629_ (.A(_12690_),
    .B(_12692_),
    .S(_12693_),
    .Z(_12694_));
 NAND2_X1 _18630_ (.A1(_11948_),
    .A2(_12694_),
    .ZN(_12695_));
 NAND2_X1 _18631_ (.A1(_11953_),
    .A2(_00816_),
    .ZN(_12696_));
 OAI21_X1 _18632_ (.A(_12696_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .B2(_12037_),
    .ZN(_12697_));
 OAI221_X1 _18633_ (.A(_12200_),
    .B1(_00815_),
    .B2(_10716_),
    .C1(_12697_),
    .C2(_11942_),
    .ZN(_12698_));
 AND3_X1 _18634_ (.A1(_10436_),
    .A2(_12695_),
    .A3(_12698_),
    .ZN(_12699_));
 MUX2_X1 _18635_ (.A(_00825_),
    .B(_00827_),
    .S(_12628_),
    .Z(_12700_));
 MUX2_X1 _18636_ (.A(_00826_),
    .B(_00828_),
    .S(_12628_),
    .Z(_12701_));
 MUX2_X1 _18637_ (.A(_12700_),
    .B(_12701_),
    .S(_12630_),
    .Z(_12702_));
 MUX2_X1 _18638_ (.A(_00817_),
    .B(_00819_),
    .S(_12628_),
    .Z(_12703_));
 BUF_X4 _18639_ (.A(net393),
    .Z(_12704_));
 MUX2_X1 _18640_ (.A(_00818_),
    .B(_00820_),
    .S(_12704_),
    .Z(_12705_));
 MUX2_X1 _18641_ (.A(_12703_),
    .B(_12705_),
    .S(_12630_),
    .Z(_12706_));
 MUX2_X1 _18642_ (.A(_12702_),
    .B(_12706_),
    .S(_11931_),
    .Z(_12707_));
 NOR2_X1 _18643_ (.A1(_12449_),
    .A2(_12707_),
    .ZN(_12708_));
 NOR3_X2 _18644_ (.A1(_11928_),
    .A2(_12699_),
    .A3(_12708_),
    .ZN(_12709_));
 MUX2_X1 _18645_ (.A(_00837_),
    .B(_00839_),
    .S(_11962_),
    .Z(_12710_));
 MUX2_X1 _18646_ (.A(_00838_),
    .B(_00840_),
    .S(_11938_),
    .Z(_12711_));
 MUX2_X1 _18647_ (.A(_12710_),
    .B(_12711_),
    .S(_11964_),
    .Z(_12712_));
 MUX2_X1 _18648_ (.A(_00829_),
    .B(_00831_),
    .S(_11962_),
    .Z(_12713_));
 MUX2_X1 _18649_ (.A(_00830_),
    .B(_00832_),
    .S(_11938_),
    .Z(_12714_));
 MUX2_X1 _18650_ (.A(_12713_),
    .B(_12714_),
    .S(_12693_),
    .Z(_12715_));
 MUX2_X1 _18651_ (.A(_12712_),
    .B(_12715_),
    .S(_11969_),
    .Z(_12716_));
 MUX2_X1 _18652_ (.A(_00841_),
    .B(_00843_),
    .S(_11938_),
    .Z(_12717_));
 MUX2_X1 _18653_ (.A(_00842_),
    .B(_00844_),
    .S(_12689_),
    .Z(_12718_));
 MUX2_X1 _18654_ (.A(_12717_),
    .B(_12718_),
    .S(_12693_),
    .Z(_12719_));
 MUX2_X1 _18655_ (.A(_00833_),
    .B(_00835_),
    .S(_12689_),
    .Z(_12720_));
 MUX2_X1 _18656_ (.A(_00834_),
    .B(_00836_),
    .S(_12691_),
    .Z(_12721_));
 MUX2_X1 _18657_ (.A(_12720_),
    .B(_12721_),
    .S(_12693_),
    .Z(_12722_));
 MUX2_X1 _18658_ (.A(_12719_),
    .B(_12722_),
    .S(_11969_),
    .Z(_12723_));
 MUX2_X1 _18659_ (.A(_12716_),
    .B(_12723_),
    .S(_12649_),
    .Z(_12724_));
 AOI21_X4 _18660_ (.A(_12709_),
    .B1(_12724_),
    .B2(_11929_),
    .ZN(_12725_));
 OAI21_X1 _18661_ (.A(_11922_),
    .B1(_11995_),
    .B2(_12725_),
    .ZN(_12726_));
 NOR2_X2 _18662_ (.A1(_12688_),
    .A2(_12726_),
    .ZN(_16008_));
 MUX2_X1 _18663_ (.A(_00821_),
    .B(_00823_),
    .S(_11597_),
    .Z(_12727_));
 MUX2_X1 _18664_ (.A(_00822_),
    .B(_00824_),
    .S(_11597_),
    .Z(_12728_));
 MUX2_X1 _18665_ (.A(_12727_),
    .B(_12728_),
    .S(_10788_),
    .Z(_12729_));
 AOI21_X1 _18666_ (.A(_10831_),
    .B1(_12729_),
    .B2(_11533_),
    .ZN(_12730_));
 NAND2_X1 _18667_ (.A1(_10602_),
    .A2(_00816_),
    .ZN(_12731_));
 OAI21_X1 _18668_ (.A(_12731_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .B2(_10622_),
    .ZN(_12732_));
 OAI22_X1 _18669_ (.A1(_00815_),
    .A2(_10758_),
    .B1(_12732_),
    .B2(_10581_),
    .ZN(_12733_));
 OAI21_X1 _18670_ (.A(_12730_),
    .B1(_12733_),
    .B2(_11533_),
    .ZN(_12734_));
 MUX2_X1 _18671_ (.A(_00837_),
    .B(_00839_),
    .S(_11546_),
    .Z(_12735_));
 MUX2_X1 _18672_ (.A(_00838_),
    .B(_00840_),
    .S(_11546_),
    .Z(_12736_));
 MUX2_X1 _18673_ (.A(_12735_),
    .B(_12736_),
    .S(_10595_),
    .Z(_12737_));
 MUX2_X1 _18674_ (.A(_00829_),
    .B(_00831_),
    .S(_11546_),
    .Z(_12738_));
 MUX2_X1 _18675_ (.A(_00830_),
    .B(_00832_),
    .S(_11546_),
    .Z(_12739_));
 MUX2_X1 _18676_ (.A(_12738_),
    .B(_12739_),
    .S(_10595_),
    .Z(_12740_));
 MUX2_X1 _18677_ (.A(_12737_),
    .B(_12740_),
    .S(_11358_),
    .Z(_12741_));
 MUX2_X1 _18678_ (.A(_00841_),
    .B(_00843_),
    .S(_11642_),
    .Z(_12742_));
 MUX2_X1 _18679_ (.A(_00842_),
    .B(_00844_),
    .S(_11642_),
    .Z(_12743_));
 MUX2_X1 _18680_ (.A(_12742_),
    .B(_12743_),
    .S(_10862_),
    .Z(_12744_));
 MUX2_X1 _18681_ (.A(_00833_),
    .B(_00835_),
    .S(_11642_),
    .Z(_12745_));
 MUX2_X1 _18682_ (.A(_00834_),
    .B(_00836_),
    .S(_10858_),
    .Z(_12746_));
 MUX2_X1 _18683_ (.A(_12745_),
    .B(_12746_),
    .S(_10862_),
    .Z(_12747_));
 MUX2_X1 _18684_ (.A(_12744_),
    .B(_12747_),
    .S(_11357_),
    .Z(_12748_));
 MUX2_X1 _18685_ (.A(_00825_),
    .B(_00827_),
    .S(_10858_),
    .Z(_12749_));
 MUX2_X1 _18686_ (.A(_00826_),
    .B(_00828_),
    .S(_10858_),
    .Z(_12750_));
 MUX2_X1 _18687_ (.A(_12749_),
    .B(_12750_),
    .S(_10862_),
    .Z(_12751_));
 MUX2_X1 _18688_ (.A(_00817_),
    .B(_00819_),
    .S(_10858_),
    .Z(_12752_));
 MUX2_X1 _18689_ (.A(_00818_),
    .B(_00820_),
    .S(_10858_),
    .Z(_12753_));
 MUX2_X1 _18690_ (.A(_12752_),
    .B(_12753_),
    .S(_10862_),
    .Z(_12754_));
 MUX2_X1 _18691_ (.A(_12751_),
    .B(_12754_),
    .S(_11357_),
    .Z(_12755_));
 MUX2_X1 _18692_ (.A(_12748_),
    .B(_12755_),
    .S(_10575_),
    .Z(_12756_));
 OAI221_X2 _18693_ (.A(_12734_),
    .B1(_11371_),
    .B2(_12741_),
    .C1(_12756_),
    .C2(_10609_),
    .ZN(_12757_));
 NAND2_X1 _18694_ (.A1(_11596_),
    .A2(net362),
    .ZN(_12758_));
 AND2_X1 _18695_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(_11593_),
    .ZN(_12759_));
 AOI22_X4 _18696_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(_10741_),
    .B1(_10683_),
    .B2(_12759_),
    .ZN(_12760_));
 NAND2_X4 _18697_ (.A1(_12758_),
    .A2(_12760_),
    .ZN(_16009_));
 INV_X2 _18698_ (.A(_16009_),
    .ZN(_16005_));
 BUF_X2 _18699_ (.A(_15454_),
    .Z(_12761_));
 INV_X1 _18700_ (.A(_12761_),
    .ZN(_12762_));
 INV_X1 _18701_ (.A(_15445_),
    .ZN(_12763_));
 INV_X1 _18702_ (.A(_12592_),
    .ZN(_12764_));
 OAI21_X1 _18703_ (.A(_12763_),
    .B1(_12598_),
    .B2(_12764_),
    .ZN(_12765_));
 BUF_X2 _18704_ (.A(_15450_),
    .Z(_12766_));
 AOI21_X2 _18705_ (.A(_15449_),
    .B1(_12765_),
    .B2(_12766_),
    .ZN(_12767_));
 INV_X1 _18706_ (.A(_12766_),
    .ZN(_12768_));
 NOR3_X2 _18707_ (.A1(_12594_),
    .A2(_12764_),
    .A3(_12768_),
    .ZN(_12769_));
 NAND2_X1 _18708_ (.A1(_12429_),
    .A2(_12769_),
    .ZN(_12770_));
 OAI21_X1 _18709_ (.A(_12767_),
    .B1(_12770_),
    .B2(_12437_),
    .ZN(_12771_));
 XNOR2_X2 _18710_ (.A(_12771_),
    .B(_12762_),
    .ZN(\alu_adder_result_ex[21] ));
 NAND2_X1 _18711_ (.A1(_12595_),
    .A2(_12608_),
    .ZN(_12772_));
 AOI21_X4 _18712_ (.A(_15445_),
    .B1(_15441_),
    .B2(_12592_),
    .ZN(_12773_));
 INV_X1 _18713_ (.A(_12773_),
    .ZN(_12774_));
 NOR3_X1 _18714_ (.A1(_12766_),
    .A2(_12772_),
    .A3(_12774_),
    .ZN(_12775_));
 AND3_X2 _18715_ (.A1(_12603_),
    .A2(_12605_),
    .A3(_12775_),
    .ZN(_12776_));
 INV_X1 _18716_ (.A(_12769_),
    .ZN(_12777_));
 AOI21_X4 _18717_ (.A(_12777_),
    .B1(_12605_),
    .B2(_12603_),
    .ZN(_12778_));
 AOI21_X1 _18718_ (.A(_12766_),
    .B1(_12592_),
    .B2(_12593_),
    .ZN(_12779_));
 NAND2_X1 _18719_ (.A1(_12773_),
    .A2(_12779_),
    .ZN(_12780_));
 OAI221_X2 _18720_ (.A(_12780_),
    .B1(_12777_),
    .B2(_12609_),
    .C1(_12768_),
    .C2(_12773_),
    .ZN(_12781_));
 NOR3_X4 _18721_ (.A1(_12776_),
    .A2(_12778_),
    .A3(_12781_),
    .ZN(\alu_adder_result_ex[20] ));
 AOI21_X1 _18722_ (.A(_12613_),
    .B1(_12614_),
    .B2(_11989_),
    .ZN(_12782_));
 MUX2_X1 _18723_ (.A(_00852_),
    .B(_00854_),
    .S(_12112_),
    .Z(_12783_));
 NOR2_X1 _18724_ (.A1(_11956_),
    .A2(_12783_),
    .ZN(_12784_));
 MUX2_X1 _18725_ (.A(_00853_),
    .B(_00855_),
    .S(_12112_),
    .Z(_12785_));
 NOR2_X1 _18726_ (.A1(_10697_),
    .A2(_12785_),
    .ZN(_12786_));
 NOR3_X1 _18727_ (.A1(_11932_),
    .A2(_12784_),
    .A3(_12786_),
    .ZN(_12787_));
 INV_X1 _18728_ (.A(_00846_),
    .ZN(_12788_));
 NOR2_X1 _18729_ (.A1(_11978_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .ZN(_12789_));
 AOI21_X1 _18730_ (.A(_12789_),
    .B1(_00847_),
    .B2(_11939_),
    .ZN(_12790_));
 AOI221_X1 _18731_ (.A(_10468_),
    .B1(_12788_),
    .B2(_11949_),
    .C1(_12790_),
    .C2(_12207_),
    .ZN(_12791_));
 NOR3_X1 _18732_ (.A1(_12649_),
    .A2(_12787_),
    .A3(_12791_),
    .ZN(_12792_));
 MUX2_X1 _18733_ (.A(_00856_),
    .B(_00858_),
    .S(_12111_),
    .Z(_12793_));
 BUF_X4 _18734_ (.A(net393),
    .Z(_12794_));
 MUX2_X1 _18735_ (.A(_00857_),
    .B(_00859_),
    .S(_12794_),
    .Z(_12795_));
 BUF_X4 _18736_ (.A(_10466_),
    .Z(_12796_));
 MUX2_X1 _18737_ (.A(_12793_),
    .B(_12795_),
    .S(_12796_),
    .Z(_12797_));
 MUX2_X1 _18738_ (.A(_00848_),
    .B(_00850_),
    .S(_12794_),
    .Z(_12798_));
 MUX2_X1 _18739_ (.A(_00849_),
    .B(_00851_),
    .S(_11943_),
    .Z(_12799_));
 MUX2_X1 _18740_ (.A(_12798_),
    .B(_12799_),
    .S(_12796_),
    .Z(_12800_));
 MUX2_X1 _18741_ (.A(_12797_),
    .B(_12800_),
    .S(_12124_),
    .Z(_12801_));
 NOR2_X1 _18742_ (.A1(_12117_),
    .A2(_12801_),
    .ZN(_12802_));
 NOR3_X2 _18743_ (.A1(_11991_),
    .A2(_12792_),
    .A3(_12802_),
    .ZN(_12803_));
 BUF_X32 _18744_ (.A(net326),
    .Z(_12804_));
 MUX2_X1 _18745_ (.A(_00868_),
    .B(_00870_),
    .S(_12804_),
    .Z(_12805_));
 BUF_X32 _18746_ (.A(net326),
    .Z(_12806_));
 MUX2_X1 _18747_ (.A(_00869_),
    .B(_00871_),
    .S(_12806_),
    .Z(_12807_));
 BUF_X4 _18748_ (.A(_11933_),
    .Z(_12808_));
 MUX2_X1 _18749_ (.A(_12805_),
    .B(_12807_),
    .S(_12808_),
    .Z(_12809_));
 MUX2_X1 _18750_ (.A(_00860_),
    .B(_00862_),
    .S(_12806_),
    .Z(_12810_));
 BUF_X32 _18751_ (.A(net326),
    .Z(_12811_));
 MUX2_X1 _18752_ (.A(_00861_),
    .B(_00863_),
    .S(_12811_),
    .Z(_12812_));
 MUX2_X1 _18753_ (.A(_12810_),
    .B(_12812_),
    .S(_12808_),
    .Z(_12813_));
 MUX2_X1 _18754_ (.A(_12809_),
    .B(_12813_),
    .S(_12017_),
    .Z(_12814_));
 MUX2_X1 _18755_ (.A(_00872_),
    .B(_00874_),
    .S(_12806_),
    .Z(_12815_));
 MUX2_X1 _18756_ (.A(_00873_),
    .B(_00875_),
    .S(_12811_),
    .Z(_12816_));
 MUX2_X1 _18757_ (.A(_12815_),
    .B(_12816_),
    .S(_12359_),
    .Z(_12817_));
 MUX2_X1 _18758_ (.A(_00864_),
    .B(_00866_),
    .S(_12811_),
    .Z(_12818_));
 MUX2_X1 _18759_ (.A(_00865_),
    .B(_00867_),
    .S(_12356_),
    .Z(_12819_));
 MUX2_X1 _18760_ (.A(_12818_),
    .B(_12819_),
    .S(_12359_),
    .Z(_12820_));
 MUX2_X1 _18761_ (.A(_12817_),
    .B(_12820_),
    .S(_12005_),
    .Z(_12821_));
 MUX2_X2 _18762_ (.A(_12814_),
    .B(_12821_),
    .S(_11930_),
    .Z(_12822_));
 AOI21_X4 _18763_ (.A(_12803_),
    .B1(_11992_),
    .B2(_12822_),
    .ZN(_12823_));
 OAI21_X1 _18764_ (.A(_11921_),
    .B1(_11994_),
    .B2(_12823_),
    .ZN(_12824_));
 NOR2_X2 _18765_ (.A1(_12782_),
    .A2(_12824_),
    .ZN(_16016_));
 NAND2_X1 _18766_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(_11632_),
    .ZN(_12825_));
 MUX2_X1 _18767_ (.A(_00872_),
    .B(_00874_),
    .S(_10585_),
    .Z(_12826_));
 MUX2_X1 _18768_ (.A(_00873_),
    .B(_00875_),
    .S(_10585_),
    .Z(_12827_));
 MUX2_X1 _18769_ (.A(_12826_),
    .B(_12827_),
    .S(_10786_),
    .Z(_12828_));
 MUX2_X1 _18770_ (.A(_00864_),
    .B(_00866_),
    .S(_10585_),
    .Z(_12829_));
 MUX2_X1 _18771_ (.A(_00865_),
    .B(_00867_),
    .S(_10585_),
    .Z(_12830_));
 MUX2_X1 _18772_ (.A(_12829_),
    .B(_12830_),
    .S(_10786_),
    .Z(_12831_));
 MUX2_X1 _18773_ (.A(_12828_),
    .B(_12831_),
    .S(_10827_),
    .Z(_12832_));
 NAND2_X1 _18774_ (.A1(_11676_),
    .A2(_12832_),
    .ZN(_12833_));
 MUX2_X1 _18775_ (.A(_00868_),
    .B(_00870_),
    .S(_11545_),
    .Z(_12834_));
 MUX2_X1 _18776_ (.A(_00869_),
    .B(_00871_),
    .S(_11545_),
    .Z(_12835_));
 MUX2_X1 _18777_ (.A(_12834_),
    .B(_12835_),
    .S(_10594_),
    .Z(_12836_));
 MUX2_X1 _18778_ (.A(_00860_),
    .B(_00861_),
    .S(_10843_),
    .Z(_12837_));
 MUX2_X1 _18779_ (.A(_00862_),
    .B(_00863_),
    .S(_10795_),
    .Z(_12838_));
 AOI222_X2 _18780_ (.A1(_10643_),
    .A2(_12836_),
    .B1(_12837_),
    .B2(_10785_),
    .C1(_12838_),
    .C2(_10794_),
    .ZN(_12839_));
 AOI21_X4 _18781_ (.A(_10783_),
    .B1(_12833_),
    .B2(_12839_),
    .ZN(_12840_));
 MUX2_X1 _18782_ (.A(_00852_),
    .B(_00854_),
    .S(_11362_),
    .Z(_12841_));
 NOR2_X1 _18783_ (.A1(_11534_),
    .A2(_12841_),
    .ZN(_12842_));
 MUX2_X1 _18784_ (.A(_00853_),
    .B(_00855_),
    .S(_11362_),
    .Z(_12843_));
 NOR2_X1 _18785_ (.A1(_10579_),
    .A2(_12843_),
    .ZN(_12844_));
 NOR3_X1 _18786_ (.A1(_11357_),
    .A2(_12842_),
    .A3(_12844_),
    .ZN(_12845_));
 NOR2_X1 _18787_ (.A1(_10612_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .ZN(_12846_));
 AOI21_X1 _18788_ (.A(_12846_),
    .B1(_00847_),
    .B2(_11771_),
    .ZN(_12847_));
 AOI221_X2 _18789_ (.A(_10765_),
    .B1(_12788_),
    .B2(_10822_),
    .C1(_12847_),
    .C2(_10795_),
    .ZN(_12848_));
 NOR3_X2 _18790_ (.A1(_10751_),
    .A2(_12845_),
    .A3(_12848_),
    .ZN(_12849_));
 MUX2_X1 _18791_ (.A(_00856_),
    .B(_00858_),
    .S(_11778_),
    .Z(_12850_));
 MUX2_X1 _18792_ (.A(_00857_),
    .B(_00859_),
    .S(_11778_),
    .Z(_12851_));
 MUX2_X1 _18793_ (.A(_12850_),
    .B(_12851_),
    .S(_10839_),
    .Z(_12852_));
 MUX2_X1 _18794_ (.A(_00848_),
    .B(_00850_),
    .S(_11778_),
    .Z(_12853_));
 MUX2_X1 _18795_ (.A(_00849_),
    .B(_00851_),
    .S(_11778_),
    .Z(_12854_));
 MUX2_X1 _18796_ (.A(_12853_),
    .B(_12854_),
    .S(_10861_),
    .Z(_12855_));
 MUX2_X1 _18797_ (.A(_12852_),
    .B(_12855_),
    .S(_11662_),
    .Z(_12856_));
 NOR2_X2 _18798_ (.A1(_11775_),
    .A2(_12856_),
    .ZN(_12857_));
 NOR3_X4 _18799_ (.A1(_11370_),
    .A2(_12849_),
    .A3(_12857_),
    .ZN(_12858_));
 OR2_X4 _18800_ (.A1(_12840_),
    .A2(_12858_),
    .ZN(_12859_));
 NAND2_X1 _18801_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(_10564_),
    .ZN(_12860_));
 OAI221_X2 _18802_ (.A(_12825_),
    .B1(_12859_),
    .B2(_10814_),
    .C1(_12860_),
    .C2(_10747_),
    .ZN(_16017_));
 INV_X2 _18803_ (.A(_16017_),
    .ZN(_16013_));
 AOI21_X1 _18804_ (.A(_12613_),
    .B1(_12614_),
    .B2(_12041_),
    .ZN(_12861_));
 MUX2_X1 _18805_ (.A(_00883_),
    .B(_00885_),
    .S(_12112_),
    .Z(_12862_));
 NOR2_X1 _18806_ (.A1(_11956_),
    .A2(_12862_),
    .ZN(_12863_));
 MUX2_X1 _18807_ (.A(_00884_),
    .B(_00886_),
    .S(_12112_),
    .Z(_12864_));
 NOR2_X1 _18808_ (.A1(_10697_),
    .A2(_12864_),
    .ZN(_12865_));
 NOR3_X1 _18809_ (.A1(_11932_),
    .A2(_12863_),
    .A3(_12865_),
    .ZN(_12866_));
 INV_X1 _18810_ (.A(_00877_),
    .ZN(_12867_));
 NOR2_X1 _18811_ (.A1(_11978_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .ZN(_12868_));
 AOI21_X1 _18812_ (.A(_12868_),
    .B1(_00878_),
    .B2(_11939_),
    .ZN(_12869_));
 AOI221_X2 _18813_ (.A(_10468_),
    .B1(_12867_),
    .B2(_11949_),
    .C1(_12869_),
    .C2(_12207_),
    .ZN(_12870_));
 NOR3_X1 _18814_ (.A1(_12649_),
    .A2(_12866_),
    .A3(_12870_),
    .ZN(_12871_));
 MUX2_X1 _18815_ (.A(_00887_),
    .B(_00889_),
    .S(_12111_),
    .Z(_12872_));
 MUX2_X1 _18816_ (.A(_00888_),
    .B(_00890_),
    .S(_12794_),
    .Z(_12873_));
 MUX2_X1 _18817_ (.A(_12872_),
    .B(_12873_),
    .S(_12796_),
    .Z(_12874_));
 MUX2_X1 _18818_ (.A(_00879_),
    .B(_00881_),
    .S(_12794_),
    .Z(_12875_));
 MUX2_X1 _18819_ (.A(_00880_),
    .B(_00882_),
    .S(_12794_),
    .Z(_12876_));
 MUX2_X1 _18820_ (.A(_12875_),
    .B(_12876_),
    .S(_12796_),
    .Z(_12877_));
 MUX2_X1 _18821_ (.A(_12874_),
    .B(_12877_),
    .S(_12124_),
    .Z(_12878_));
 NOR2_X1 _18822_ (.A1(_12117_),
    .A2(_12878_),
    .ZN(_12879_));
 NOR3_X2 _18823_ (.A1(_11991_),
    .A2(_12871_),
    .A3(_12879_),
    .ZN(_12880_));
 MUX2_X1 _18824_ (.A(_00899_),
    .B(_00901_),
    .S(net429),
    .Z(_12881_));
 MUX2_X1 _18825_ (.A(_00900_),
    .B(_00902_),
    .S(_12806_),
    .Z(_12882_));
 MUX2_X1 _18826_ (.A(_12881_),
    .B(_12882_),
    .S(_12808_),
    .Z(_12883_));
 MUX2_X1 _18827_ (.A(_00891_),
    .B(_00893_),
    .S(_12804_),
    .Z(_12884_));
 MUX2_X1 _18828_ (.A(_00892_),
    .B(_00894_),
    .S(net435),
    .Z(_12885_));
 MUX2_X1 _18829_ (.A(_12884_),
    .B(_12885_),
    .S(_12808_),
    .Z(_12886_));
 MUX2_X1 _18830_ (.A(_12883_),
    .B(_12886_),
    .S(_12017_),
    .Z(_12887_));
 MUX2_X1 _18831_ (.A(_00903_),
    .B(_00905_),
    .S(_12806_),
    .Z(_12888_));
 MUX2_X1 _18832_ (.A(_00904_),
    .B(_00906_),
    .S(_12811_),
    .Z(_12889_));
 MUX2_X1 _18833_ (.A(_12888_),
    .B(_12889_),
    .S(_12359_),
    .Z(_12890_));
 MUX2_X1 _18834_ (.A(_00895_),
    .B(_00897_),
    .S(net435),
    .Z(_12891_));
 MUX2_X1 _18835_ (.A(_00896_),
    .B(_00898_),
    .S(_12356_),
    .Z(_12892_));
 MUX2_X1 _18836_ (.A(_12891_),
    .B(_12892_),
    .S(_12359_),
    .Z(_12893_));
 MUX2_X1 _18837_ (.A(_12890_),
    .B(_12893_),
    .S(_12005_),
    .Z(_12894_));
 MUX2_X2 _18838_ (.A(_12887_),
    .B(_12894_),
    .S(_11930_),
    .Z(_12895_));
 AOI21_X4 _18839_ (.A(_12880_),
    .B1(_12895_),
    .B2(_11992_),
    .ZN(_12896_));
 OAI21_X1 _18840_ (.A(_11921_),
    .B1(_11994_),
    .B2(_12896_),
    .ZN(_12897_));
 NOR2_X2 _18841_ (.A1(_12861_),
    .A2(_12897_),
    .ZN(_16021_));
 NAND2_X1 _18842_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(_11632_),
    .ZN(_12898_));
 MUX2_X1 _18843_ (.A(_00899_),
    .B(_00901_),
    .S(_11641_),
    .Z(_12899_));
 MUX2_X1 _18844_ (.A(_00900_),
    .B(_00902_),
    .S(_11641_),
    .Z(_12900_));
 MUX2_X1 _18845_ (.A(_12899_),
    .B(_12900_),
    .S(_10861_),
    .Z(_12901_));
 MUX2_X1 _18846_ (.A(_00891_),
    .B(_00893_),
    .S(_10857_),
    .Z(_12902_));
 MUX2_X1 _18847_ (.A(_00892_),
    .B(_00894_),
    .S(_10857_),
    .Z(_12903_));
 MUX2_X1 _18848_ (.A(_12902_),
    .B(_12903_),
    .S(_10593_),
    .Z(_12904_));
 MUX2_X1 _18849_ (.A(_12901_),
    .B(_12904_),
    .S(_10568_),
    .Z(_12905_));
 NOR2_X1 _18850_ (.A1(_10751_),
    .A2(_12905_),
    .ZN(_12906_));
 MUX2_X1 _18851_ (.A(_00903_),
    .B(_00905_),
    .S(_11778_),
    .Z(_12907_));
 MUX2_X1 _18852_ (.A(_00904_),
    .B(_00906_),
    .S(_11641_),
    .Z(_12908_));
 MUX2_X1 _18853_ (.A(_12907_),
    .B(_12908_),
    .S(_10861_),
    .Z(_12909_));
 MUX2_X1 _18854_ (.A(_00895_),
    .B(_00897_),
    .S(_11641_),
    .Z(_12910_));
 MUX2_X1 _18855_ (.A(_00896_),
    .B(_00898_),
    .S(_11641_),
    .Z(_12911_));
 MUX2_X1 _18856_ (.A(_12910_),
    .B(_12911_),
    .S(_10861_),
    .Z(_12912_));
 MUX2_X1 _18857_ (.A(_12909_),
    .B(_12912_),
    .S(_11662_),
    .Z(_12913_));
 NOR2_X1 _18858_ (.A1(_11775_),
    .A2(_12913_),
    .ZN(_12914_));
 NOR3_X4 _18859_ (.A1(_10783_),
    .A2(_12906_),
    .A3(_12914_),
    .ZN(_12915_));
 MUX2_X1 _18860_ (.A(_00883_),
    .B(_00885_),
    .S(_11362_),
    .Z(_12916_));
 NOR2_X1 _18861_ (.A1(_11534_),
    .A2(_12916_),
    .ZN(_12917_));
 MUX2_X1 _18862_ (.A(_00884_),
    .B(_00886_),
    .S(_12498_),
    .Z(_12918_));
 NOR2_X1 _18863_ (.A1(_10579_),
    .A2(_12918_),
    .ZN(_12919_));
 NOR3_X1 _18864_ (.A1(_10827_),
    .A2(_12917_),
    .A3(_12919_),
    .ZN(_12920_));
 NOR2_X1 _18865_ (.A1(_11567_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .ZN(_12921_));
 AOI21_X1 _18866_ (.A(_12921_),
    .B1(_00878_),
    .B2(_11771_),
    .ZN(_12922_));
 AOI221_X2 _18867_ (.A(_10764_),
    .B1(_12867_),
    .B2(_10822_),
    .C1(_12922_),
    .C2(_10786_),
    .ZN(_12923_));
 NOR3_X2 _18868_ (.A1(_10832_),
    .A2(_12920_),
    .A3(_12923_),
    .ZN(_12924_));
 MUX2_X1 _18869_ (.A(_00887_),
    .B(_00889_),
    .S(_10790_),
    .Z(_12925_));
 MUX2_X1 _18870_ (.A(_00888_),
    .B(_00890_),
    .S(_10790_),
    .Z(_12926_));
 MUX2_X1 _18871_ (.A(_12925_),
    .B(_12926_),
    .S(_10833_),
    .Z(_12927_));
 MUX2_X1 _18872_ (.A(_00879_),
    .B(_00881_),
    .S(_10790_),
    .Z(_12928_));
 MUX2_X1 _18873_ (.A(_00880_),
    .B(_00882_),
    .S(_10790_),
    .Z(_12929_));
 MUX2_X1 _18874_ (.A(_12928_),
    .B(_12929_),
    .S(_10833_),
    .Z(_12930_));
 MUX2_X1 _18875_ (.A(_12927_),
    .B(_12930_),
    .S(_11662_),
    .Z(_12931_));
 NOR2_X1 _18876_ (.A1(_11775_),
    .A2(_12931_),
    .ZN(_12932_));
 NOR3_X4 _18877_ (.A1(_11370_),
    .A2(_12924_),
    .A3(_12932_),
    .ZN(_12933_));
 OR2_X2 _18878_ (.A1(_12915_),
    .A2(_12933_),
    .ZN(_12934_));
 CLKBUF_X2 _18879_ (.A(\cs_registers_i.pc_id_i[23] ),
    .Z(_12935_));
 NAND2_X1 _18880_ (.A1(_12935_),
    .A2(_10564_),
    .ZN(_12936_));
 OAI221_X2 _18881_ (.A(_12898_),
    .B1(_12934_),
    .B2(_10814_),
    .C1(_12936_),
    .C2(_10746_),
    .ZN(_16020_));
 INV_X2 _18882_ (.A(_16020_),
    .ZN(_16024_));
 INV_X1 _18883_ (.A(_15462_),
    .ZN(_12937_));
 INV_X1 _18884_ (.A(_15457_),
    .ZN(_12938_));
 NAND4_X1 _18885_ (.A1(_12592_),
    .A2(_12766_),
    .A3(_12761_),
    .A4(_15458_),
    .ZN(_12939_));
 INV_X1 _18886_ (.A(_15449_),
    .ZN(_12940_));
 OAI21_X1 _18887_ (.A(_12940_),
    .B1(_12763_),
    .B2(_12768_),
    .ZN(_12941_));
 AOI21_X1 _18888_ (.A(_15453_),
    .B1(_12941_),
    .B2(_12761_),
    .ZN(_12942_));
 INV_X1 _18889_ (.A(_15458_),
    .ZN(_12943_));
 OAI221_X2 _18890_ (.A(_12938_),
    .B1(_12600_),
    .B2(_12939_),
    .C1(_12942_),
    .C2(_12943_),
    .ZN(_12944_));
 XNOR2_X2 _18891_ (.A(_12937_),
    .B(_12944_),
    .ZN(\alu_adder_result_ex[23] ));
 OAI21_X1 _18892_ (.A(_12940_),
    .B1(_12773_),
    .B2(_12768_),
    .ZN(_12945_));
 AOI21_X2 _18893_ (.A(_15453_),
    .B1(_12945_),
    .B2(_12761_),
    .ZN(_12946_));
 NAND2_X1 _18894_ (.A1(_12761_),
    .A2(_12769_),
    .ZN(_12947_));
 OAI21_X1 _18895_ (.A(_12946_),
    .B1(_12947_),
    .B2(_12610_),
    .ZN(_12948_));
 XNOR2_X2 _18896_ (.A(_12943_),
    .B(_12948_),
    .ZN(_12949_));
 BUF_X8 _18897_ (.A(_12949_),
    .Z(\alu_adder_result_ex[22] ));
 AOI21_X1 _18898_ (.A(_12613_),
    .B1(_12614_),
    .B2(_11992_),
    .ZN(_12950_));
 MUX2_X1 _18899_ (.A(_00914_),
    .B(_00916_),
    .S(_12112_),
    .Z(_12951_));
 NOR2_X1 _18900_ (.A1(_11956_),
    .A2(_12951_),
    .ZN(_12952_));
 MUX2_X1 _18901_ (.A(_00915_),
    .B(_00917_),
    .S(_11978_),
    .Z(_12953_));
 NOR2_X1 _18902_ (.A1(_10697_),
    .A2(_12953_),
    .ZN(_12954_));
 NOR3_X1 _18903_ (.A1(_11932_),
    .A2(_12952_),
    .A3(_12954_),
    .ZN(_12955_));
 INV_X1 _18904_ (.A(_00908_),
    .ZN(_12956_));
 NOR2_X1 _18905_ (.A1(_11978_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .ZN(_12957_));
 AOI21_X1 _18906_ (.A(_12957_),
    .B1(_00909_),
    .B2(_11939_),
    .ZN(_12958_));
 AOI221_X2 _18907_ (.A(_10468_),
    .B1(_12956_),
    .B2(_10964_),
    .C1(_12958_),
    .C2(_12207_),
    .ZN(_12959_));
 NOR3_X1 _18908_ (.A1(_12649_),
    .A2(_12955_),
    .A3(_12959_),
    .ZN(_12960_));
 MUX2_X1 _18909_ (.A(_00918_),
    .B(_00920_),
    .S(_12111_),
    .Z(_12961_));
 MUX2_X1 _18910_ (.A(_00919_),
    .B(_00921_),
    .S(_12111_),
    .Z(_12962_));
 MUX2_X1 _18911_ (.A(_12961_),
    .B(_12962_),
    .S(_12796_),
    .Z(_12963_));
 MUX2_X1 _18912_ (.A(_00910_),
    .B(_00912_),
    .S(_12111_),
    .Z(_12964_));
 MUX2_X1 _18913_ (.A(_00911_),
    .B(_00913_),
    .S(_12794_),
    .Z(_12965_));
 MUX2_X1 _18914_ (.A(_12964_),
    .B(_12965_),
    .S(_12796_),
    .Z(_12966_));
 MUX2_X1 _18915_ (.A(_12963_),
    .B(_12966_),
    .S(_12124_),
    .Z(_12967_));
 NOR2_X1 _18916_ (.A1(_12117_),
    .A2(_12967_),
    .ZN(_12968_));
 NOR3_X2 _18917_ (.A1(_11991_),
    .A2(_12960_),
    .A3(_12968_),
    .ZN(_12969_));
 MUX2_X1 _18918_ (.A(_00930_),
    .B(_00932_),
    .S(net429),
    .Z(_12970_));
 MUX2_X1 _18919_ (.A(_00931_),
    .B(_00933_),
    .S(net429),
    .Z(_12971_));
 MUX2_X1 _18920_ (.A(_12970_),
    .B(_12971_),
    .S(_12012_),
    .Z(_12972_));
 MUX2_X1 _18921_ (.A(_00922_),
    .B(_00924_),
    .S(net429),
    .Z(_12973_));
 MUX2_X1 _18922_ (.A(_00923_),
    .B(_00925_),
    .S(_12804_),
    .Z(_12974_));
 MUX2_X1 _18923_ (.A(_12973_),
    .B(_12974_),
    .S(_12012_),
    .Z(_12975_));
 MUX2_X1 _18924_ (.A(_12972_),
    .B(_12975_),
    .S(_12017_),
    .Z(_12976_));
 MUX2_X1 _18925_ (.A(_00934_),
    .B(_00936_),
    .S(_12010_),
    .Z(_12977_));
 MUX2_X1 _18926_ (.A(_00935_),
    .B(_00937_),
    .S(_12804_),
    .Z(_12978_));
 MUX2_X1 _18927_ (.A(_12977_),
    .B(_12978_),
    .S(_12808_),
    .Z(_12979_));
 MUX2_X1 _18928_ (.A(_00926_),
    .B(_00928_),
    .S(_12804_),
    .Z(_12980_));
 MUX2_X1 _18929_ (.A(_00927_),
    .B(_00929_),
    .S(_12811_),
    .Z(_12981_));
 MUX2_X1 _18930_ (.A(_12980_),
    .B(_12981_),
    .S(_12808_),
    .Z(_12982_));
 MUX2_X1 _18931_ (.A(_12979_),
    .B(_12982_),
    .S(_12017_),
    .Z(_12983_));
 MUX2_X2 _18932_ (.A(_12976_),
    .B(_12983_),
    .S(_11930_),
    .Z(_12984_));
 AOI21_X4 _18933_ (.A(_12969_),
    .B1(_12984_),
    .B2(_11929_),
    .ZN(_12985_));
 OAI21_X1 _18934_ (.A(_11921_),
    .B1(_11994_),
    .B2(_12985_),
    .ZN(_12986_));
 NOR2_X2 _18935_ (.A1(_12950_),
    .A2(_12986_),
    .ZN(_16032_));
 NAND2_X1 _18936_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(_11632_),
    .ZN(_12987_));
 MUX2_X1 _18937_ (.A(_00930_),
    .B(_00932_),
    .S(_10857_),
    .Z(_12988_));
 MUX2_X1 _18938_ (.A(_00931_),
    .B(_00933_),
    .S(_10857_),
    .Z(_12989_));
 MUX2_X1 _18939_ (.A(_12988_),
    .B(_12989_),
    .S(_10593_),
    .Z(_12990_));
 MUX2_X1 _18940_ (.A(_00922_),
    .B(_00924_),
    .S(_10857_),
    .Z(_12991_));
 MUX2_X1 _18941_ (.A(_00923_),
    .B(_00925_),
    .S(_10857_),
    .Z(_12992_));
 MUX2_X1 _18942_ (.A(_12991_),
    .B(_12992_),
    .S(_10593_),
    .Z(_12993_));
 MUX2_X1 _18943_ (.A(_12990_),
    .B(_12993_),
    .S(_10568_),
    .Z(_12994_));
 NOR2_X1 _18944_ (.A1(_10751_),
    .A2(_12994_),
    .ZN(_12995_));
 MUX2_X1 _18945_ (.A(_00934_),
    .B(_00936_),
    .S(_11641_),
    .Z(_12996_));
 MUX2_X1 _18946_ (.A(_00935_),
    .B(_00937_),
    .S(_11641_),
    .Z(_12997_));
 MUX2_X1 _18947_ (.A(_12996_),
    .B(_12997_),
    .S(_10861_),
    .Z(_12998_));
 MUX2_X1 _18948_ (.A(_00926_),
    .B(_00928_),
    .S(_11641_),
    .Z(_12999_));
 MUX2_X1 _18949_ (.A(_00927_),
    .B(_00929_),
    .S(_11641_),
    .Z(_13000_));
 MUX2_X1 _18950_ (.A(_12999_),
    .B(_13000_),
    .S(_10861_),
    .Z(_13001_));
 MUX2_X1 _18951_ (.A(_12998_),
    .B(_13001_),
    .S(_11662_),
    .Z(_13002_));
 NOR2_X1 _18952_ (.A1(_10608_),
    .A2(_13002_),
    .ZN(_13003_));
 NOR3_X4 _18953_ (.A1(_10783_),
    .A2(_12995_),
    .A3(_13003_),
    .ZN(_13004_));
 MUX2_X1 _18954_ (.A(_00914_),
    .B(_00916_),
    .S(_11362_),
    .Z(_13005_));
 NOR2_X1 _18955_ (.A1(_11534_),
    .A2(_13005_),
    .ZN(_13006_));
 MUX2_X1 _18956_ (.A(_00915_),
    .B(_00917_),
    .S(_12498_),
    .Z(_13007_));
 NOR2_X1 _18957_ (.A1(_10579_),
    .A2(_13007_),
    .ZN(_13008_));
 NOR3_X1 _18958_ (.A1(_10827_),
    .A2(_13006_),
    .A3(_13008_),
    .ZN(_13009_));
 NOR2_X1 _18959_ (.A1(_11567_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .ZN(_13010_));
 AOI21_X1 _18960_ (.A(_13010_),
    .B1(_00909_),
    .B2(_11771_),
    .ZN(_13011_));
 AOI221_X2 _18961_ (.A(_10764_),
    .B1(_12956_),
    .B2(_10822_),
    .C1(_13011_),
    .C2(_10786_),
    .ZN(_13012_));
 NOR3_X2 _18962_ (.A1(_10832_),
    .A2(_13009_),
    .A3(_13012_),
    .ZN(_13013_));
 MUX2_X1 _18963_ (.A(_00918_),
    .B(_00920_),
    .S(_10790_),
    .Z(_13014_));
 MUX2_X1 _18964_ (.A(_00919_),
    .B(_00921_),
    .S(_11776_),
    .Z(_13015_));
 MUX2_X1 _18965_ (.A(_13014_),
    .B(_13015_),
    .S(_10839_),
    .Z(_13016_));
 MUX2_X1 _18966_ (.A(_00910_),
    .B(_00912_),
    .S(_11776_),
    .Z(_13017_));
 MUX2_X1 _18967_ (.A(_00911_),
    .B(_00913_),
    .S(_11776_),
    .Z(_13018_));
 MUX2_X1 _18968_ (.A(_13017_),
    .B(_13018_),
    .S(_10839_),
    .Z(_13019_));
 MUX2_X1 _18969_ (.A(_13016_),
    .B(_13019_),
    .S(_11662_),
    .Z(_13020_));
 NOR2_X2 _18970_ (.A1(_11775_),
    .A2(_13020_),
    .ZN(_13021_));
 NOR3_X4 _18971_ (.A1(_11370_),
    .A2(_13013_),
    .A3(_13021_),
    .ZN(_13022_));
 OR2_X2 _18972_ (.A1(_13004_),
    .A2(_13022_),
    .ZN(_13023_));
 CLKBUF_X2 _18973_ (.A(\cs_registers_i.pc_id_i[24] ),
    .Z(_13024_));
 NAND2_X1 _18974_ (.A1(_13024_),
    .A2(_10564_),
    .ZN(_13025_));
 OAI221_X2 _18975_ (.A(_12987_),
    .B1(_13023_),
    .B2(_10814_),
    .C1(_13025_),
    .C2(_10747_),
    .ZN(_16033_));
 INV_X2 _18976_ (.A(_16033_),
    .ZN(_16029_));
 AOI21_X1 _18977_ (.A(_12613_),
    .B1(_12614_),
    .B2(_10873_),
    .ZN(_13026_));
 MUX2_X1 _18978_ (.A(_00945_),
    .B(_00947_),
    .S(_12112_),
    .Z(_13027_));
 NOR2_X1 _18979_ (.A1(_11956_),
    .A2(_13027_),
    .ZN(_13028_));
 MUX2_X1 _18980_ (.A(_00946_),
    .B(_00948_),
    .S(_12112_),
    .Z(_13029_));
 NOR2_X1 _18981_ (.A1(_10697_),
    .A2(_13029_),
    .ZN(_13030_));
 NOR3_X1 _18982_ (.A1(_11932_),
    .A2(_13028_),
    .A3(_13030_),
    .ZN(_13031_));
 INV_X1 _18983_ (.A(_00939_),
    .ZN(_13032_));
 NOR2_X1 _18984_ (.A1(_11978_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .ZN(_13033_));
 AOI21_X1 _18985_ (.A(_13033_),
    .B1(_00940_),
    .B2(_11939_),
    .ZN(_13034_));
 AOI221_X2 _18986_ (.A(_10468_),
    .B1(_13032_),
    .B2(_11949_),
    .C1(_13034_),
    .C2(_12207_),
    .ZN(_13035_));
 NOR3_X1 _18987_ (.A1(_12649_),
    .A2(_13031_),
    .A3(_13035_),
    .ZN(_13036_));
 MUX2_X1 _18988_ (.A(_00949_),
    .B(_00951_),
    .S(_12111_),
    .Z(_13037_));
 MUX2_X1 _18989_ (.A(_00950_),
    .B(_00952_),
    .S(_12794_),
    .Z(_13038_));
 MUX2_X1 _18990_ (.A(_13037_),
    .B(_13038_),
    .S(_12796_),
    .Z(_13039_));
 MUX2_X1 _18991_ (.A(_00941_),
    .B(_00943_),
    .S(_12794_),
    .Z(_13040_));
 MUX2_X1 _18992_ (.A(_00942_),
    .B(_00944_),
    .S(_11943_),
    .Z(_13041_));
 MUX2_X1 _18993_ (.A(_13040_),
    .B(_13041_),
    .S(_11955_),
    .Z(_13042_));
 MUX2_X1 _18994_ (.A(_13039_),
    .B(_13042_),
    .S(_12124_),
    .Z(_13043_));
 NOR2_X1 _18995_ (.A1(_12117_),
    .A2(_13043_),
    .ZN(_13044_));
 NOR3_X2 _18996_ (.A1(_11991_),
    .A2(_13036_),
    .A3(_13044_),
    .ZN(_13045_));
 MUX2_X1 _18997_ (.A(_00961_),
    .B(_00963_),
    .S(net436),
    .Z(_13046_));
 MUX2_X1 _18998_ (.A(_00962_),
    .B(_00964_),
    .S(net433),
    .Z(_13047_));
 MUX2_X1 _18999_ (.A(_13046_),
    .B(_13047_),
    .S(_12808_),
    .Z(_13048_));
 MUX2_X1 _19000_ (.A(_00953_),
    .B(_00955_),
    .S(net433),
    .Z(_13049_));
 MUX2_X1 _19001_ (.A(_00954_),
    .B(_00956_),
    .S(net435),
    .Z(_13050_));
 MUX2_X1 _19002_ (.A(_13049_),
    .B(_13050_),
    .S(_12359_),
    .Z(_13051_));
 MUX2_X1 _19003_ (.A(_13048_),
    .B(_13051_),
    .S(_12017_),
    .Z(_13052_));
 MUX2_X1 _19004_ (.A(_00965_),
    .B(_00967_),
    .S(net433),
    .Z(_13053_));
 MUX2_X1 _19005_ (.A(_00966_),
    .B(_00968_),
    .S(net402),
    .Z(_13054_));
 MUX2_X1 _19006_ (.A(_13053_),
    .B(_13054_),
    .S(_12359_),
    .Z(_13055_));
 MUX2_X1 _19007_ (.A(_00957_),
    .B(_00959_),
    .S(net402),
    .Z(_13056_));
 MUX2_X1 _19008_ (.A(_00958_),
    .B(_00960_),
    .S(net402),
    .Z(_13057_));
 MUX2_X1 _19009_ (.A(_13056_),
    .B(_13057_),
    .S(_12359_),
    .Z(_13058_));
 MUX2_X1 _19010_ (.A(_13055_),
    .B(_13058_),
    .S(_12005_),
    .Z(_13059_));
 MUX2_X2 _19011_ (.A(_13052_),
    .B(_13059_),
    .S(_11930_),
    .Z(_13060_));
 AOI21_X4 _19012_ (.A(_13045_),
    .B1(_11992_),
    .B2(_13060_),
    .ZN(_13061_));
 OAI21_X1 _19013_ (.A(_11921_),
    .B1(_11994_),
    .B2(_13061_),
    .ZN(_13062_));
 NOR2_X2 _19014_ (.A1(_13026_),
    .A2(_13062_),
    .ZN(_16037_));
 AND3_X1 _19015_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(_10563_),
    .A3(_10682_),
    .ZN(_13063_));
 MUX2_X1 _19016_ (.A(_00965_),
    .B(_00967_),
    .S(_11385_),
    .Z(_13064_));
 MUX2_X1 _19017_ (.A(_00966_),
    .B(_00968_),
    .S(_11385_),
    .Z(_13065_));
 MUX2_X1 _19018_ (.A(_13064_),
    .B(_13065_),
    .S(_11383_),
    .Z(_13066_));
 MUX2_X1 _19019_ (.A(_00957_),
    .B(_00959_),
    .S(_11385_),
    .Z(_13067_));
 MUX2_X1 _19020_ (.A(_00958_),
    .B(_00960_),
    .S(_11385_),
    .Z(_13068_));
 MUX2_X1 _19021_ (.A(_13067_),
    .B(_13068_),
    .S(_11383_),
    .Z(_13069_));
 MUX2_X1 _19022_ (.A(_13066_),
    .B(_13069_),
    .S(_10568_),
    .Z(_13070_));
 NAND2_X1 _19023_ (.A1(_11676_),
    .A2(_13070_),
    .ZN(_13071_));
 MUX2_X1 _19024_ (.A(_00961_),
    .B(_00963_),
    .S(_11362_),
    .Z(_13072_));
 MUX2_X1 _19025_ (.A(_00962_),
    .B(_00964_),
    .S(_11362_),
    .Z(_13073_));
 MUX2_X1 _19026_ (.A(_13072_),
    .B(_13073_),
    .S(_10839_),
    .Z(_13074_));
 MUX2_X1 _19027_ (.A(_00955_),
    .B(_00956_),
    .S(_10795_),
    .Z(_13075_));
 MUX2_X1 _19028_ (.A(_00953_),
    .B(_00954_),
    .S(_10786_),
    .Z(_13076_));
 AOI222_X2 _19029_ (.A1(_10643_),
    .A2(_13074_),
    .B1(_13075_),
    .B2(_10794_),
    .C1(_13076_),
    .C2(_10785_),
    .ZN(_13077_));
 AOI21_X4 _19030_ (.A(_10575_),
    .B1(_13071_),
    .B2(_13077_),
    .ZN(_13078_));
 MUX2_X1 _19031_ (.A(_00945_),
    .B(_00947_),
    .S(_12498_),
    .Z(_13079_));
 NOR2_X1 _19032_ (.A1(_10594_),
    .A2(_13079_),
    .ZN(_13080_));
 MUX2_X1 _19033_ (.A(_00946_),
    .B(_00948_),
    .S(_11567_),
    .Z(_13081_));
 NOR2_X1 _19034_ (.A1(_10579_),
    .A2(_13081_),
    .ZN(_13082_));
 NOR3_X1 _19035_ (.A1(_10827_),
    .A2(_13080_),
    .A3(_13082_),
    .ZN(_13083_));
 NOR2_X1 _19036_ (.A1(_10618_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .ZN(_13084_));
 AOI21_X1 _19037_ (.A(_13084_),
    .B1(_00940_),
    .B2(_11545_),
    .ZN(_13085_));
 AOI221_X2 _19038_ (.A(_10764_),
    .B1(_13032_),
    .B2(_10821_),
    .C1(_13085_),
    .C2(_10626_),
    .ZN(_13086_));
 NOR3_X2 _19039_ (.A1(_10832_),
    .A2(_13083_),
    .A3(_13086_),
    .ZN(_13087_));
 MUX2_X1 _19040_ (.A(_00949_),
    .B(_00951_),
    .S(_11655_),
    .Z(_13088_));
 MUX2_X1 _19041_ (.A(_00950_),
    .B(_00952_),
    .S(_11655_),
    .Z(_13089_));
 MUX2_X1 _19042_ (.A(_13088_),
    .B(_13089_),
    .S(_10833_),
    .Z(_13090_));
 MUX2_X1 _19043_ (.A(_00941_),
    .B(_00943_),
    .S(_11655_),
    .Z(_13091_));
 MUX2_X1 _19044_ (.A(_00942_),
    .B(_00944_),
    .S(_11655_),
    .Z(_13092_));
 MUX2_X1 _19045_ (.A(_13091_),
    .B(_13092_),
    .S(_10833_),
    .Z(_13093_));
 MUX2_X1 _19046_ (.A(_13090_),
    .B(_13093_),
    .S(_10567_),
    .Z(_13094_));
 NOR2_X2 _19047_ (.A1(_11775_),
    .A2(_13094_),
    .ZN(_13095_));
 NOR3_X4 _19048_ (.A1(_11370_),
    .A2(_13087_),
    .A3(_13095_),
    .ZN(_13096_));
 NOR2_X4 _19049_ (.A1(_13078_),
    .A2(_13096_),
    .ZN(_13097_));
 AOI221_X2 _19050_ (.A(_13063_),
    .B1(_13097_),
    .B2(_10816_),
    .C1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .C2(_11632_),
    .ZN(_13098_));
 BUF_X4 _19051_ (.A(_13098_),
    .Z(_16040_));
 CLKBUF_X2 _19052_ (.A(_15470_),
    .Z(_13099_));
 INV_X1 _19053_ (.A(_15461_),
    .ZN(_13100_));
 AOI21_X1 _19054_ (.A(_15457_),
    .B1(_15453_),
    .B2(_15458_),
    .ZN(_13101_));
 OAI21_X1 _19055_ (.A(_13100_),
    .B1(_13101_),
    .B2(_12937_),
    .ZN(_13102_));
 CLKBUF_X2 _19056_ (.A(_15466_),
    .Z(_13103_));
 AOI21_X2 _19057_ (.A(_15465_),
    .B1(_13102_),
    .B2(_13103_),
    .ZN(_13104_));
 NAND2_X1 _19058_ (.A1(_15458_),
    .A2(_15462_),
    .ZN(_13105_));
 NOR2_X1 _19059_ (.A1(_12762_),
    .A2(_13105_),
    .ZN(_13106_));
 AND3_X1 _19060_ (.A1(_13103_),
    .A2(_12769_),
    .A3(_13106_),
    .ZN(_13107_));
 NAND2_X1 _19061_ (.A1(_12429_),
    .A2(_13107_),
    .ZN(_13108_));
 NAND2_X1 _19062_ (.A1(_13103_),
    .A2(_13106_),
    .ZN(_13109_));
 OAI221_X2 _19063_ (.A(_13104_),
    .B1(_13108_),
    .B2(_12437_),
    .C1(_12767_),
    .C2(_13109_),
    .ZN(_13110_));
 XNOR2_X2 _19064_ (.A(_13110_),
    .B(_13099_),
    .ZN(_13111_));
 INV_X4 _19065_ (.A(_13111_),
    .ZN(\alu_adder_result_ex[25] ));
 AOI21_X1 _19066_ (.A(_15453_),
    .B1(_15449_),
    .B2(_12761_),
    .ZN(_13112_));
 OAI21_X1 _19067_ (.A(_12938_),
    .B1(_13112_),
    .B2(_12943_),
    .ZN(_13113_));
 AOI21_X1 _19068_ (.A(_15461_),
    .B1(_13113_),
    .B2(_15462_),
    .ZN(_13114_));
 NAND2_X1 _19069_ (.A1(_12766_),
    .A2(_13106_),
    .ZN(_13115_));
 AOI21_X1 _19070_ (.A(_12774_),
    .B1(_12592_),
    .B2(_12593_),
    .ZN(_13116_));
 OAI21_X1 _19071_ (.A(_13114_),
    .B1(_13115_),
    .B2(_13116_),
    .ZN(_13117_));
 NAND2_X1 _19072_ (.A1(_12773_),
    .A2(_13114_),
    .ZN(_13118_));
 NAND3_X1 _19073_ (.A1(_12603_),
    .A2(_12605_),
    .A3(_12609_),
    .ZN(_13119_));
 OAI21_X2 _19074_ (.A(_13117_),
    .B1(_13118_),
    .B2(_13119_),
    .ZN(_13120_));
 XNOR2_X2 _19075_ (.A(_13103_),
    .B(_13120_),
    .ZN(_13121_));
 BUF_X4 _19076_ (.A(_13121_),
    .Z(\alu_adder_result_ex[24] ));
 AOI21_X1 _19077_ (.A(_12613_),
    .B1(_12614_),
    .B2(_10874_),
    .ZN(_13122_));
 MUX2_X1 _19078_ (.A(_00976_),
    .B(_00978_),
    .S(net436),
    .Z(_13123_));
 MUX2_X1 _19079_ (.A(_00977_),
    .B(_00979_),
    .S(net433),
    .Z(_13124_));
 MUX2_X1 _19080_ (.A(_13123_),
    .B(_13124_),
    .S(_12808_),
    .Z(_13125_));
 NAND2_X1 _19081_ (.A1(_12041_),
    .A2(_13125_),
    .ZN(_13126_));
 NAND2_X1 _19082_ (.A1(_11953_),
    .A2(_00971_),
    .ZN(_13127_));
 OAI21_X1 _19083_ (.A(_13127_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B2(_12034_),
    .ZN(_13128_));
 OAI221_X1 _19084_ (.A(_12200_),
    .B1(_00970_),
    .B2(_10716_),
    .C1(_13128_),
    .C2(_11942_),
    .ZN(_13129_));
 AND3_X1 _19085_ (.A1(_12449_),
    .A2(_13126_),
    .A3(_13129_),
    .ZN(_13130_));
 MUX2_X1 _19086_ (.A(_00980_),
    .B(_00982_),
    .S(_12111_),
    .Z(_13131_));
 MUX2_X1 _19087_ (.A(_00981_),
    .B(_00983_),
    .S(_12111_),
    .Z(_13132_));
 MUX2_X1 _19088_ (.A(_13131_),
    .B(_13132_),
    .S(_12796_),
    .Z(_13133_));
 MUX2_X1 _19089_ (.A(_00972_),
    .B(_00974_),
    .S(_12794_),
    .Z(_13134_));
 MUX2_X1 _19090_ (.A(_00973_),
    .B(_00975_),
    .S(_12794_),
    .Z(_13135_));
 MUX2_X1 _19091_ (.A(_13134_),
    .B(_13135_),
    .S(_12796_),
    .Z(_13136_));
 MUX2_X1 _19092_ (.A(_13133_),
    .B(_13136_),
    .S(_12124_),
    .Z(_13137_));
 NOR2_X1 _19093_ (.A1(_12117_),
    .A2(_13137_),
    .ZN(_13138_));
 NOR3_X2 _19094_ (.A1(_11991_),
    .A2(_13130_),
    .A3(_13138_),
    .ZN(_13139_));
 MUX2_X1 _19095_ (.A(_00992_),
    .B(_00994_),
    .S(net429),
    .Z(_13140_));
 MUX2_X1 _19096_ (.A(_00993_),
    .B(_00995_),
    .S(net436),
    .Z(_13141_));
 MUX2_X1 _19097_ (.A(_13140_),
    .B(_13141_),
    .S(_12012_),
    .Z(_13142_));
 MUX2_X1 _19098_ (.A(_00984_),
    .B(_00986_),
    .S(net436),
    .Z(_13143_));
 MUX2_X1 _19099_ (.A(_00985_),
    .B(_00987_),
    .S(net433),
    .Z(_13144_));
 MUX2_X1 _19100_ (.A(_13143_),
    .B(_13144_),
    .S(_12808_),
    .Z(_13145_));
 MUX2_X1 _19101_ (.A(_13142_),
    .B(_13145_),
    .S(_12017_),
    .Z(_13146_));
 MUX2_X1 _19102_ (.A(_00996_),
    .B(_00998_),
    .S(net436),
    .Z(_13147_));
 MUX2_X1 _19103_ (.A(_00997_),
    .B(_00999_),
    .S(net435),
    .Z(_13148_));
 MUX2_X1 _19104_ (.A(_13147_),
    .B(_13148_),
    .S(_12808_),
    .Z(_13149_));
 MUX2_X1 _19105_ (.A(_00988_),
    .B(_00990_),
    .S(net435),
    .Z(_13150_));
 MUX2_X1 _19106_ (.A(_00989_),
    .B(_00991_),
    .S(net402),
    .Z(_13151_));
 MUX2_X1 _19107_ (.A(_13150_),
    .B(_13151_),
    .S(_12359_),
    .Z(_13152_));
 MUX2_X1 _19108_ (.A(_13149_),
    .B(_13152_),
    .S(_12005_),
    .Z(_13153_));
 MUX2_X2 _19109_ (.A(_13146_),
    .B(_13153_),
    .S(_11930_),
    .Z(_13154_));
 AOI21_X4 _19110_ (.A(_13139_),
    .B1(_11929_),
    .B2(_13154_),
    .ZN(_13155_));
 OAI21_X1 _19111_ (.A(_11921_),
    .B1(_11994_),
    .B2(_13155_),
    .ZN(_13156_));
 NOR2_X2 _19112_ (.A1(_13122_),
    .A2(_13156_),
    .ZN(_16048_));
 MUX2_X1 _19113_ (.A(_00976_),
    .B(_00978_),
    .S(_10600_),
    .Z(_13157_));
 MUX2_X1 _19114_ (.A(_00977_),
    .B(_00979_),
    .S(_10600_),
    .Z(_13158_));
 MUX2_X1 _19115_ (.A(_13157_),
    .B(_13158_),
    .S(_10628_),
    .Z(_13159_));
 AOI21_X1 _19116_ (.A(_10831_),
    .B1(_13159_),
    .B2(_10766_),
    .ZN(_13160_));
 NAND2_X1 _19117_ (.A1(_10615_),
    .A2(_00971_),
    .ZN(_13161_));
 OAI21_X1 _19118_ (.A(_13161_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B2(_10602_),
    .ZN(_13162_));
 OAI22_X1 _19119_ (.A1(_00970_),
    .A2(_10757_),
    .B1(_13162_),
    .B2(_10581_),
    .ZN(_13163_));
 OAI21_X1 _19120_ (.A(_13160_),
    .B1(_13163_),
    .B2(_11533_),
    .ZN(_13164_));
 MUX2_X1 _19121_ (.A(_00992_),
    .B(_00994_),
    .S(_10613_),
    .Z(_13165_));
 MUX2_X1 _19122_ (.A(_00993_),
    .B(_00995_),
    .S(_10613_),
    .Z(_13166_));
 MUX2_X1 _19123_ (.A(_13165_),
    .B(_13166_),
    .S(_11877_),
    .Z(_13167_));
 MUX2_X1 _19124_ (.A(_00984_),
    .B(_00986_),
    .S(_10613_),
    .Z(_13168_));
 MUX2_X1 _19125_ (.A(_00985_),
    .B(_00987_),
    .S(_10613_),
    .Z(_13169_));
 MUX2_X1 _19126_ (.A(_13168_),
    .B(_13169_),
    .S(_11877_),
    .Z(_13170_));
 MUX2_X2 _19127_ (.A(_13167_),
    .B(_13170_),
    .S(_10828_),
    .Z(_13171_));
 MUX2_X1 _19128_ (.A(_00996_),
    .B(_00998_),
    .S(_10612_),
    .Z(_13172_));
 MUX2_X1 _19129_ (.A(_00997_),
    .B(_00999_),
    .S(_10612_),
    .Z(_13173_));
 MUX2_X1 _19130_ (.A(_13172_),
    .B(_13173_),
    .S(_10843_),
    .Z(_13174_));
 MUX2_X1 _19131_ (.A(_00988_),
    .B(_00990_),
    .S(_10612_),
    .Z(_13175_));
 MUX2_X1 _19132_ (.A(_00989_),
    .B(_00991_),
    .S(_10612_),
    .Z(_13176_));
 MUX2_X1 _19133_ (.A(_13175_),
    .B(_13176_),
    .S(_10843_),
    .Z(_13177_));
 MUX2_X1 _19134_ (.A(_13174_),
    .B(_13177_),
    .S(_11357_),
    .Z(_13178_));
 MUX2_X1 _19135_ (.A(_00980_),
    .B(_00982_),
    .S(_10612_),
    .Z(_13179_));
 MUX2_X1 _19136_ (.A(_00981_),
    .B(_00983_),
    .S(_10612_),
    .Z(_13180_));
 MUX2_X1 _19137_ (.A(_13179_),
    .B(_13180_),
    .S(_10843_),
    .Z(_13181_));
 MUX2_X1 _19138_ (.A(_00972_),
    .B(_00974_),
    .S(_10612_),
    .Z(_13182_));
 MUX2_X1 _19139_ (.A(_00973_),
    .B(_00975_),
    .S(_10612_),
    .Z(_13183_));
 MUX2_X1 _19140_ (.A(_13182_),
    .B(_13183_),
    .S(_10843_),
    .Z(_13184_));
 MUX2_X1 _19141_ (.A(_13181_),
    .B(_13184_),
    .S(_11357_),
    .Z(_13185_));
 MUX2_X1 _19142_ (.A(_13178_),
    .B(_13185_),
    .S(_10575_),
    .Z(_13186_));
 OAI221_X2 _19143_ (.A(_13164_),
    .B1(_13171_),
    .B2(_11371_),
    .C1(_10609_),
    .C2(_13186_),
    .ZN(_13187_));
 AND2_X1 _19144_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(_11593_),
    .ZN(_13188_));
 AOI222_X4 _19145_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(_10397_),
    .B1(_11596_),
    .B2(net351),
    .C1(_13188_),
    .C2(_10870_),
    .ZN(_16045_));
 AOI21_X1 _19146_ (.A(_12613_),
    .B1(_12614_),
    .B2(_10500_),
    .ZN(_13189_));
 BUF_X4 _19147_ (.A(net437),
    .Z(_13190_));
 MUX2_X1 _19148_ (.A(_01007_),
    .B(_01009_),
    .S(_13190_),
    .Z(_13191_));
 MUX2_X1 _19149_ (.A(_01008_),
    .B(_01010_),
    .S(_12008_),
    .Z(_13192_));
 BUF_X4 _19150_ (.A(_11933_),
    .Z(_13193_));
 MUX2_X1 _19151_ (.A(_13191_),
    .B(_13192_),
    .S(_13193_),
    .Z(_13194_));
 NAND2_X1 _19152_ (.A1(_12041_),
    .A2(_13194_),
    .ZN(_13195_));
 NAND2_X1 _19153_ (.A1(_11953_),
    .A2(_01002_),
    .ZN(_13196_));
 OAI21_X1 _19154_ (.A(_13196_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .B2(_12034_),
    .ZN(_13197_));
 OAI221_X1 _19155_ (.A(_12200_),
    .B1(_01001_),
    .B2(_10716_),
    .C1(_13197_),
    .C2(_11942_),
    .ZN(_13198_));
 AND3_X1 _19156_ (.A1(_12449_),
    .A2(_13195_),
    .A3(_13198_),
    .ZN(_13199_));
 MUX2_X1 _19157_ (.A(_01011_),
    .B(_01013_),
    .S(_12628_),
    .Z(_13200_));
 MUX2_X1 _19158_ (.A(_01012_),
    .B(_01014_),
    .S(_12704_),
    .Z(_13201_));
 MUX2_X1 _19159_ (.A(_13200_),
    .B(_13201_),
    .S(_12630_),
    .Z(_13202_));
 MUX2_X1 _19160_ (.A(_01003_),
    .B(_01005_),
    .S(_12704_),
    .Z(_13203_));
 MUX2_X1 _19161_ (.A(_01004_),
    .B(_01006_),
    .S(_12111_),
    .Z(_13204_));
 MUX2_X1 _19162_ (.A(_13203_),
    .B(_13204_),
    .S(_12796_),
    .Z(_13205_));
 MUX2_X1 _19163_ (.A(_13202_),
    .B(_13205_),
    .S(_12124_),
    .Z(_13206_));
 NOR2_X1 _19164_ (.A1(_12117_),
    .A2(_13206_),
    .ZN(_13207_));
 NOR3_X2 _19165_ (.A1(_11928_),
    .A2(_13199_),
    .A3(_13207_),
    .ZN(_13208_));
 MUX2_X1 _19166_ (.A(_01023_),
    .B(_01025_),
    .S(net428),
    .Z(_13209_));
 MUX2_X1 _19167_ (.A(_01024_),
    .B(_01026_),
    .S(net434),
    .Z(_13210_));
 MUX2_X1 _19168_ (.A(_13209_),
    .B(_13210_),
    .S(_12693_),
    .Z(_13211_));
 MUX2_X1 _19169_ (.A(_01015_),
    .B(_01017_),
    .S(_12691_),
    .Z(_13212_));
 MUX2_X1 _19170_ (.A(_01016_),
    .B(_01018_),
    .S(_13190_),
    .Z(_13213_));
 MUX2_X1 _19171_ (.A(_13212_),
    .B(_13213_),
    .S(_13193_),
    .Z(_13214_));
 MUX2_X1 _19172_ (.A(_13211_),
    .B(_13214_),
    .S(_11969_),
    .Z(_13215_));
 MUX2_X1 _19173_ (.A(_01027_),
    .B(_01029_),
    .S(_12691_),
    .Z(_13216_));
 MUX2_X1 _19174_ (.A(_01028_),
    .B(_01030_),
    .S(_13190_),
    .Z(_13217_));
 MUX2_X1 _19175_ (.A(_13216_),
    .B(_13217_),
    .S(_13193_),
    .Z(_13218_));
 MUX2_X1 _19176_ (.A(_01019_),
    .B(_01021_),
    .S(_13190_),
    .Z(_13219_));
 MUX2_X1 _19177_ (.A(_01020_),
    .B(_01022_),
    .S(_12008_),
    .Z(_13220_));
 MUX2_X1 _19178_ (.A(_13219_),
    .B(_13220_),
    .S(_12012_),
    .Z(_13221_));
 MUX2_X1 _19179_ (.A(_13218_),
    .B(_13221_),
    .S(_12017_),
    .Z(_13222_));
 MUX2_X1 _19180_ (.A(_13215_),
    .B(_13222_),
    .S(_12649_),
    .Z(_13223_));
 AOI21_X4 _19181_ (.A(_13208_),
    .B1(_11929_),
    .B2(_13223_),
    .ZN(_13224_));
 OAI21_X1 _19182_ (.A(_11921_),
    .B1(_11994_),
    .B2(_13224_),
    .ZN(_13225_));
 NOR2_X2 _19183_ (.A1(_13189_),
    .A2(_13225_),
    .ZN(_16053_));
 AND2_X1 _19184_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_10564_),
    .ZN(_13226_));
 AOI22_X4 _19185_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(_10397_),
    .B1(_10683_),
    .B2(_13226_),
    .ZN(_13227_));
 NAND2_X1 _19186_ (.A1(_10622_),
    .A2(_01002_),
    .ZN(_13228_));
 OAI21_X1 _19187_ (.A(_13228_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .B2(_10616_),
    .ZN(_13229_));
 OAI221_X1 _19188_ (.A(_10576_),
    .B1(_01001_),
    .B2(_10758_),
    .C1(_13229_),
    .C2(_10582_),
    .ZN(_13230_));
 MUX2_X1 _19189_ (.A(_01015_),
    .B(_01017_),
    .S(_11547_),
    .Z(_13231_));
 MUX2_X1 _19190_ (.A(_01016_),
    .B(_01018_),
    .S(_11547_),
    .Z(_13232_));
 MUX2_X1 _19191_ (.A(_13231_),
    .B(_13232_),
    .S(_10596_),
    .Z(_13233_));
 AOI21_X1 _19192_ (.A(_11437_),
    .B1(_13233_),
    .B2(_10749_),
    .ZN(_13234_));
 NAND2_X1 _19193_ (.A1(_13230_),
    .A2(_13234_),
    .ZN(_13235_));
 MUX2_X1 _19194_ (.A(_01023_),
    .B(_01025_),
    .S(_10587_),
    .Z(_13236_));
 MUX2_X1 _19195_ (.A(_01024_),
    .B(_01026_),
    .S(_10587_),
    .Z(_13237_));
 MUX2_X1 _19196_ (.A(_13236_),
    .B(_13237_),
    .S(_10788_),
    .Z(_13238_));
 MUX2_X1 _19197_ (.A(_01007_),
    .B(_01009_),
    .S(_10620_),
    .Z(_13239_));
 MUX2_X1 _19198_ (.A(_01008_),
    .B(_01010_),
    .S(_10620_),
    .Z(_13240_));
 MUX2_X1 _19199_ (.A(_13239_),
    .B(_13240_),
    .S(_10788_),
    .Z(_13241_));
 MUX2_X1 _19200_ (.A(_13238_),
    .B(_13241_),
    .S(_10783_),
    .Z(_13242_));
 MUX2_X1 _19201_ (.A(_01027_),
    .B(_01029_),
    .S(_10585_),
    .Z(_13243_));
 MUX2_X1 _19202_ (.A(_01028_),
    .B(_01030_),
    .S(_10585_),
    .Z(_13244_));
 MUX2_X1 _19203_ (.A(_13243_),
    .B(_13244_),
    .S(_10787_),
    .Z(_13245_));
 MUX2_X1 _19204_ (.A(_01011_),
    .B(_01013_),
    .S(_10585_),
    .Z(_13246_));
 MUX2_X1 _19205_ (.A(_01012_),
    .B(_01014_),
    .S(_10585_),
    .Z(_13247_));
 MUX2_X1 _19206_ (.A(_13246_),
    .B(_13247_),
    .S(_10787_),
    .Z(_13248_));
 MUX2_X1 _19207_ (.A(_13245_),
    .B(_13248_),
    .S(_10574_),
    .Z(_13249_));
 MUX2_X1 _19208_ (.A(_01019_),
    .B(_01021_),
    .S(_10585_),
    .Z(_13250_));
 MUX2_X1 _19209_ (.A(_01020_),
    .B(_01022_),
    .S(_10585_),
    .Z(_13251_));
 MUX2_X1 _19210_ (.A(_13250_),
    .B(_13251_),
    .S(_10787_),
    .Z(_13252_));
 MUX2_X1 _19211_ (.A(_01003_),
    .B(_01005_),
    .S(_10585_),
    .Z(_13253_));
 MUX2_X1 _19212_ (.A(_01004_),
    .B(_01006_),
    .S(_10619_),
    .Z(_13254_));
 MUX2_X1 _19213_ (.A(_13253_),
    .B(_13254_),
    .S(_10787_),
    .Z(_13255_));
 MUX2_X1 _19214_ (.A(_13252_),
    .B(_13255_),
    .S(_10574_),
    .Z(_13256_));
 MUX2_X1 _19215_ (.A(_13249_),
    .B(_13256_),
    .S(_10570_),
    .Z(_13257_));
 OAI221_X2 _19216_ (.A(_13235_),
    .B1(_11453_),
    .B2(_13242_),
    .C1(_13257_),
    .C2(_10610_),
    .ZN(_13258_));
 INV_X2 _19217_ (.A(net341),
    .ZN(_13259_));
 OAI21_X4 _19218_ (.A(_13227_),
    .B1(_13259_),
    .B2(_10814_),
    .ZN(_16052_));
 INV_X2 _19219_ (.A(_16052_),
    .ZN(_16056_));
 INV_X2 _19220_ (.A(_15478_),
    .ZN(_13260_));
 OAI21_X1 _19221_ (.A(_13104_),
    .B1(_13109_),
    .B2(_12767_),
    .ZN(_13261_));
 CLKBUF_X3 _19222_ (.A(_15474_),
    .Z(_13262_));
 AND2_X1 _19223_ (.A1(_13099_),
    .A2(_13262_),
    .ZN(_13263_));
 AOI221_X2 _19224_ (.A(_15473_),
    .B1(_13261_),
    .B2(_13263_),
    .C1(_15469_),
    .C2(_13262_),
    .ZN(_13264_));
 NAND3_X2 _19225_ (.A1(_12429_),
    .A2(_13107_),
    .A3(_13263_),
    .ZN(_13265_));
 OAI21_X4 _19226_ (.A(_13264_),
    .B1(_12437_),
    .B2(_13265_),
    .ZN(_13266_));
 XNOR2_X2 _19227_ (.A(_13266_),
    .B(_13260_),
    .ZN(\alu_adder_result_ex[27] ));
 AND2_X1 _19228_ (.A1(_13099_),
    .A2(_13107_),
    .ZN(_13267_));
 NAND2_X1 _19229_ (.A1(_13262_),
    .A2(_13267_),
    .ZN(_13268_));
 NOR2_X1 _19230_ (.A1(_12609_),
    .A2(_13268_),
    .ZN(_13269_));
 NOR2_X1 _19231_ (.A1(_13262_),
    .A2(_13267_),
    .ZN(_13270_));
 AOI21_X1 _19232_ (.A(_15469_),
    .B1(_15465_),
    .B2(_13099_),
    .ZN(_13271_));
 INV_X1 _19233_ (.A(_13271_),
    .ZN(_13272_));
 AND2_X1 _19234_ (.A1(_13103_),
    .A2(_13099_),
    .ZN(_13273_));
 OAI221_X2 _19235_ (.A(_13100_),
    .B1(_12946_),
    .B2(_13105_),
    .C1(_12938_),
    .C2(_12937_),
    .ZN(_13274_));
 AOI21_X2 _19236_ (.A(_13272_),
    .B1(_13273_),
    .B2(_13274_),
    .ZN(_13275_));
 MUX2_X1 _19237_ (.A(_13262_),
    .B(_13270_),
    .S(_13275_),
    .Z(_13276_));
 AOI21_X2 _19238_ (.A(_13268_),
    .B1(_12605_),
    .B2(_12603_),
    .ZN(_13277_));
 INV_X1 _19239_ (.A(_13262_),
    .ZN(_13278_));
 AND2_X1 _19240_ (.A1(_13278_),
    .A2(_13275_),
    .ZN(_13279_));
 AND4_X1 _19241_ (.A1(_12603_),
    .A2(_12605_),
    .A3(_12609_),
    .A4(_13279_),
    .ZN(_13280_));
 NOR4_X4 _19242_ (.A1(_13269_),
    .A2(_13280_),
    .A3(_13277_),
    .A4(_13276_),
    .ZN(\alu_adder_result_ex[26] ));
 AOI21_X1 _19243_ (.A(_12613_),
    .B1(_12614_),
    .B2(_10501_),
    .ZN(_13281_));
 MUX2_X1 _19244_ (.A(_01038_),
    .B(_01040_),
    .S(net434),
    .Z(_13282_));
 MUX2_X1 _19245_ (.A(_01039_),
    .B(_01041_),
    .S(_12008_),
    .Z(_13283_));
 MUX2_X1 _19246_ (.A(_13282_),
    .B(_13283_),
    .S(_13193_),
    .Z(_13284_));
 NAND2_X1 _19247_ (.A1(_12041_),
    .A2(_13284_),
    .ZN(_13285_));
 NAND2_X1 _19248_ (.A1(_11953_),
    .A2(_01033_),
    .ZN(_13286_));
 OAI21_X1 _19249_ (.A(_13286_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .B2(_12034_),
    .ZN(_13287_));
 OAI221_X1 _19250_ (.A(_12200_),
    .B1(_01032_),
    .B2(_10716_),
    .C1(_13287_),
    .C2(_11942_),
    .ZN(_13288_));
 AND3_X1 _19251_ (.A1(_12449_),
    .A2(_13285_),
    .A3(_13288_),
    .ZN(_13289_));
 MUX2_X1 _19252_ (.A(_01042_),
    .B(_01044_),
    .S(_12628_),
    .Z(_13290_));
 MUX2_X1 _19253_ (.A(_01043_),
    .B(_01045_),
    .S(_12704_),
    .Z(_13291_));
 MUX2_X1 _19254_ (.A(_13290_),
    .B(_13291_),
    .S(_12630_),
    .Z(_13292_));
 MUX2_X1 _19255_ (.A(_01034_),
    .B(_01036_),
    .S(_12704_),
    .Z(_13293_));
 MUX2_X1 _19256_ (.A(_01035_),
    .B(_01037_),
    .S(_12704_),
    .Z(_13294_));
 MUX2_X1 _19257_ (.A(_13293_),
    .B(_13294_),
    .S(_12630_),
    .Z(_13295_));
 MUX2_X1 _19258_ (.A(_13292_),
    .B(_13295_),
    .S(_12124_),
    .Z(_13296_));
 NOR2_X1 _19259_ (.A1(_12449_),
    .A2(_13296_),
    .ZN(_13297_));
 NOR3_X2 _19260_ (.A1(_11928_),
    .A2(_13289_),
    .A3(_13297_),
    .ZN(_13298_));
 MUX2_X1 _19261_ (.A(_01054_),
    .B(_01056_),
    .S(net428),
    .Z(_13299_));
 MUX2_X1 _19262_ (.A(_01055_),
    .B(_01057_),
    .S(net427),
    .Z(_13300_));
 MUX2_X1 _19263_ (.A(_13299_),
    .B(_13300_),
    .S(_12693_),
    .Z(_13301_));
 MUX2_X1 _19264_ (.A(_01046_),
    .B(_01048_),
    .S(net427),
    .Z(_13302_));
 MUX2_X1 _19265_ (.A(_01047_),
    .B(_01049_),
    .S(_13190_),
    .Z(_13303_));
 MUX2_X1 _19266_ (.A(_13302_),
    .B(_13303_),
    .S(_13193_),
    .Z(_13304_));
 MUX2_X1 _19267_ (.A(_13301_),
    .B(_13304_),
    .S(_11969_),
    .Z(_13305_));
 MUX2_X1 _19268_ (.A(_01058_),
    .B(_01060_),
    .S(net434),
    .Z(_13306_));
 MUX2_X1 _19269_ (.A(_01059_),
    .B(_01061_),
    .S(_13190_),
    .Z(_13307_));
 MUX2_X1 _19270_ (.A(_13306_),
    .B(_13307_),
    .S(_13193_),
    .Z(_13308_));
 MUX2_X1 _19271_ (.A(_01050_),
    .B(_01052_),
    .S(_13190_),
    .Z(_13309_));
 MUX2_X1 _19272_ (.A(_01051_),
    .B(_01053_),
    .S(_12008_),
    .Z(_13310_));
 MUX2_X1 _19273_ (.A(_13309_),
    .B(_13310_),
    .S(_12012_),
    .Z(_13311_));
 MUX2_X1 _19274_ (.A(_13308_),
    .B(_13311_),
    .S(_12017_),
    .Z(_13312_));
 MUX2_X2 _19275_ (.A(_13305_),
    .B(_13312_),
    .S(_12649_),
    .Z(_13313_));
 AOI21_X4 _19276_ (.A(_13298_),
    .B1(_11929_),
    .B2(_13313_),
    .ZN(_13314_));
 OAI21_X1 _19277_ (.A(_11921_),
    .B1(_11994_),
    .B2(_13314_),
    .ZN(_03093_));
 NOR2_X2 _19278_ (.A1(_13281_),
    .A2(_03093_),
    .ZN(_16061_));
 NAND2_X1 _19279_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(_10397_),
    .ZN(_03094_));
 MUX2_X1 _19280_ (.A(_01038_),
    .B(_01040_),
    .S(_10601_),
    .Z(_03095_));
 MUX2_X1 _19281_ (.A(_01039_),
    .B(_01041_),
    .S(_10601_),
    .Z(_03096_));
 MUX2_X1 _19282_ (.A(_03095_),
    .B(_03096_),
    .S(_10596_),
    .Z(_03097_));
 NAND2_X1 _19283_ (.A1(_10767_),
    .A2(_03097_),
    .ZN(_03098_));
 NAND2_X1 _19284_ (.A1(_10622_),
    .A2(_01033_),
    .ZN(_03099_));
 OAI21_X1 _19285_ (.A(_03099_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .B2(_10616_),
    .ZN(_03100_));
 OAI221_X2 _19286_ (.A(_10571_),
    .B1(_01032_),
    .B2(_10758_),
    .C1(_03100_),
    .C2(_10581_),
    .ZN(_03101_));
 NAND3_X2 _19287_ (.A1(_10610_),
    .A2(_03098_),
    .A3(_03101_),
    .ZN(_03102_));
 MUX2_X1 _19288_ (.A(_01042_),
    .B(_01044_),
    .S(_11547_),
    .Z(_03103_));
 MUX2_X1 _19289_ (.A(_01043_),
    .B(_01045_),
    .S(_11547_),
    .Z(_03104_));
 MUX2_X1 _19290_ (.A(_03103_),
    .B(_03104_),
    .S(_10596_),
    .Z(_03105_));
 NAND2_X1 _19291_ (.A1(_11533_),
    .A2(_03105_),
    .ZN(_03106_));
 MUX2_X1 _19292_ (.A(_01034_),
    .B(_01036_),
    .S(_11547_),
    .Z(_03107_));
 MUX2_X1 _19293_ (.A(_01035_),
    .B(_01037_),
    .S(_11547_),
    .Z(_03108_));
 MUX2_X1 _19294_ (.A(_03107_),
    .B(_03108_),
    .S(_10596_),
    .Z(_03109_));
 NAND2_X1 _19295_ (.A1(_10571_),
    .A2(_03109_),
    .ZN(_03110_));
 NAND3_X2 _19296_ (.A1(_10752_),
    .A2(_03106_),
    .A3(_03110_),
    .ZN(_03111_));
 AOI21_X4 _19297_ (.A(_10750_),
    .B1(_03102_),
    .B2(_03111_),
    .ZN(_03112_));
 MUX2_X1 _19298_ (.A(_01050_),
    .B(_01052_),
    .S(_10587_),
    .Z(_03113_));
 MUX2_X1 _19299_ (.A(_01051_),
    .B(_01053_),
    .S(_10587_),
    .Z(_03114_));
 MUX2_X1 _19300_ (.A(_03113_),
    .B(_03114_),
    .S(_10628_),
    .Z(_03115_));
 MUX2_X1 _19301_ (.A(_01048_),
    .B(_01049_),
    .S(_11535_),
    .Z(_03116_));
 MUX2_X1 _19302_ (.A(_01046_),
    .B(_01047_),
    .S(_11366_),
    .Z(_03117_));
 AOI222_X2 _19303_ (.A1(_10778_),
    .A2(_03115_),
    .B1(_03116_),
    .B2(_10794_),
    .C1(_03117_),
    .C2(_10785_),
    .ZN(_03118_));
 NAND2_X1 _19304_ (.A1(_10749_),
    .A2(_03118_),
    .ZN(_03119_));
 MUX2_X1 _19305_ (.A(_01060_),
    .B(_01061_),
    .S(_11534_),
    .Z(_03120_));
 AOI21_X2 _19306_ (.A(_11775_),
    .B1(_03120_),
    .B2(_10602_),
    .ZN(_03121_));
 MUX2_X1 _19307_ (.A(_01056_),
    .B(_01057_),
    .S(_10862_),
    .Z(_03122_));
 AOI21_X2 _19308_ (.A(_10606_),
    .B1(_03122_),
    .B2(_10621_),
    .ZN(_03123_));
 OAI21_X2 _19309_ (.A(_10759_),
    .B1(_03121_),
    .B2(_03123_),
    .ZN(_03124_));
 MUX2_X1 _19310_ (.A(_01054_),
    .B(_01055_),
    .S(_10627_),
    .Z(_03125_));
 INV_X1 _19311_ (.A(_03125_),
    .ZN(_03126_));
 MUX2_X1 _19312_ (.A(_01058_),
    .B(_01059_),
    .S(_11366_),
    .Z(_03127_));
 INV_X1 _19313_ (.A(_03127_),
    .ZN(_03128_));
 AOI221_X2 _19314_ (.A(_10570_),
    .B1(_03123_),
    .B2(_03126_),
    .C1(_03128_),
    .C2(_03121_),
    .ZN(_03129_));
 AOI21_X4 _19315_ (.A(_03119_),
    .B1(_03124_),
    .B2(_03129_),
    .ZN(_03130_));
 NOR2_X4 _19316_ (.A1(_03112_),
    .A2(_03130_),
    .ZN(_03131_));
 NAND2_X1 _19317_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_10565_),
    .ZN(_03132_));
 OAI221_X2 _19318_ (.A(_03094_),
    .B1(_03131_),
    .B2(_10814_),
    .C1(_03132_),
    .C2(_10747_),
    .ZN(_16060_));
 INV_X2 _19319_ (.A(_16060_),
    .ZN(_16064_));
 AOI21_X1 _19320_ (.A(_12613_),
    .B1(_12614_),
    .B2(_10502_),
    .ZN(_03133_));
 MUX2_X1 _19321_ (.A(_01069_),
    .B(_01071_),
    .S(net434),
    .Z(_03134_));
 MUX2_X1 _19322_ (.A(_01070_),
    .B(_01072_),
    .S(_12008_),
    .Z(_03135_));
 MUX2_X1 _19323_ (.A(_03134_),
    .B(_03135_),
    .S(_13193_),
    .Z(_03136_));
 NAND2_X1 _19324_ (.A1(_11948_),
    .A2(_03136_),
    .ZN(_03137_));
 NAND2_X1 _19325_ (.A1(_11953_),
    .A2(_01064_),
    .ZN(_03138_));
 OAI21_X1 _19326_ (.A(_03138_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .B2(_12034_),
    .ZN(_03139_));
 OAI221_X1 _19327_ (.A(_12200_),
    .B1(_01063_),
    .B2(_10716_),
    .C1(_03139_),
    .C2(_11942_),
    .ZN(_03140_));
 AND3_X1 _19328_ (.A1(_12449_),
    .A2(_03137_),
    .A3(_03140_),
    .ZN(_03141_));
 MUX2_X1 _19329_ (.A(_01073_),
    .B(_01075_),
    .S(_12628_),
    .Z(_03142_));
 MUX2_X1 _19330_ (.A(_01074_),
    .B(_01076_),
    .S(_12704_),
    .Z(_03143_));
 MUX2_X1 _19331_ (.A(_03142_),
    .B(_03143_),
    .S(_12630_),
    .Z(_03144_));
 MUX2_X1 _19332_ (.A(_01065_),
    .B(_01067_),
    .S(_12704_),
    .Z(_03145_));
 MUX2_X1 _19333_ (.A(_01066_),
    .B(_01068_),
    .S(_12704_),
    .Z(_03146_));
 MUX2_X1 _19334_ (.A(_03145_),
    .B(_03146_),
    .S(_12630_),
    .Z(_03147_));
 MUX2_X1 _19335_ (.A(_03144_),
    .B(_03147_),
    .S(_12124_),
    .Z(_03148_));
 NOR2_X1 _19336_ (.A1(_12449_),
    .A2(_03148_),
    .ZN(_03149_));
 NOR3_X2 _19337_ (.A1(_11928_),
    .A2(_03141_),
    .A3(_03149_),
    .ZN(_03150_));
 MUX2_X1 _19338_ (.A(_01085_),
    .B(_01087_),
    .S(net428),
    .Z(_03151_));
 MUX2_X1 _19339_ (.A(_01086_),
    .B(_01088_),
    .S(net427),
    .Z(_03152_));
 MUX2_X1 _19340_ (.A(_03151_),
    .B(_03152_),
    .S(_12693_),
    .Z(_03153_));
 MUX2_X1 _19341_ (.A(_01077_),
    .B(_01079_),
    .S(net427),
    .Z(_03154_));
 MUX2_X1 _19342_ (.A(_01078_),
    .B(_01080_),
    .S(_13190_),
    .Z(_03155_));
 MUX2_X1 _19343_ (.A(_03154_),
    .B(_03155_),
    .S(_13193_),
    .Z(_03156_));
 MUX2_X1 _19344_ (.A(_03153_),
    .B(_03156_),
    .S(_11969_),
    .Z(_03157_));
 MUX2_X1 _19345_ (.A(_01089_),
    .B(_01091_),
    .S(net434),
    .Z(_03158_));
 MUX2_X1 _19346_ (.A(_01090_),
    .B(_01092_),
    .S(_13190_),
    .Z(_03159_));
 MUX2_X1 _19347_ (.A(_03158_),
    .B(_03159_),
    .S(_13193_),
    .Z(_03160_));
 MUX2_X1 _19348_ (.A(_01081_),
    .B(_01083_),
    .S(_13190_),
    .Z(_03161_));
 MUX2_X1 _19349_ (.A(_01082_),
    .B(_01084_),
    .S(_12008_),
    .Z(_03162_));
 MUX2_X1 _19350_ (.A(_03161_),
    .B(_03162_),
    .S(_12012_),
    .Z(_03163_));
 MUX2_X1 _19351_ (.A(_03160_),
    .B(_03163_),
    .S(_11969_),
    .Z(_03164_));
 MUX2_X1 _19352_ (.A(_03157_),
    .B(_03164_),
    .S(_12649_),
    .Z(_03165_));
 AOI21_X4 _19353_ (.A(_03150_),
    .B1(_03165_),
    .B2(_11929_),
    .ZN(_03166_));
 OAI21_X1 _19354_ (.A(_11921_),
    .B1(_11994_),
    .B2(_03166_),
    .ZN(_03167_));
 NOR2_X2 _19355_ (.A1(_03133_),
    .A2(_03167_),
    .ZN(_16069_));
 MUX2_X1 _19356_ (.A(_01069_),
    .B(_01071_),
    .S(_10602_),
    .Z(_03168_));
 MUX2_X1 _19357_ (.A(_01070_),
    .B(_01072_),
    .S(_10602_),
    .Z(_03169_));
 MUX2_X1 _19358_ (.A(_03168_),
    .B(_03169_),
    .S(_10597_),
    .Z(_03170_));
 NAND2_X1 _19359_ (.A1(_10767_),
    .A2(_03170_),
    .ZN(_03171_));
 NAND2_X1 _19360_ (.A1(_10759_),
    .A2(_01064_),
    .ZN(_03172_));
 OAI21_X1 _19361_ (.A(_03172_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .B2(_10759_),
    .ZN(_03173_));
 OAI221_X2 _19362_ (.A(_10571_),
    .B1(_01063_),
    .B2(_10758_),
    .C1(_03173_),
    .C2(_10582_),
    .ZN(_03174_));
 NAND3_X2 _19363_ (.A1(_10610_),
    .A2(_03171_),
    .A3(_03174_),
    .ZN(_03175_));
 MUX2_X1 _19364_ (.A(_01073_),
    .B(_01075_),
    .S(_10615_),
    .Z(_03176_));
 MUX2_X1 _19365_ (.A(_01074_),
    .B(_01076_),
    .S(_10615_),
    .Z(_03177_));
 MUX2_X1 _19366_ (.A(_03176_),
    .B(_03177_),
    .S(_10597_),
    .Z(_03178_));
 NAND2_X1 _19367_ (.A1(_10767_),
    .A2(_03178_),
    .ZN(_03179_));
 MUX2_X1 _19368_ (.A(_01065_),
    .B(_01067_),
    .S(_10615_),
    .Z(_03180_));
 MUX2_X1 _19369_ (.A(_01066_),
    .B(_01068_),
    .S(_10615_),
    .Z(_03181_));
 MUX2_X1 _19370_ (.A(_03180_),
    .B(_03181_),
    .S(_10629_),
    .Z(_03182_));
 NAND2_X1 _19371_ (.A1(_10571_),
    .A2(_03182_),
    .ZN(_03183_));
 NAND3_X2 _19372_ (.A1(_10752_),
    .A2(_03179_),
    .A3(_03183_),
    .ZN(_03184_));
 AOI21_X4 _19373_ (.A(_10750_),
    .B1(_03175_),
    .B2(_03184_),
    .ZN(_03185_));
 MUX2_X1 _19374_ (.A(_01081_),
    .B(_01083_),
    .S(_10588_),
    .Z(_03186_));
 MUX2_X1 _19375_ (.A(_01082_),
    .B(_01084_),
    .S(_10588_),
    .Z(_03187_));
 MUX2_X1 _19376_ (.A(_03186_),
    .B(_03187_),
    .S(_10629_),
    .Z(_03188_));
 MUX2_X1 _19377_ (.A(_01079_),
    .B(_01080_),
    .S(_10596_),
    .Z(_03189_));
 MUX2_X1 _19378_ (.A(_01077_),
    .B(_01078_),
    .S(_10797_),
    .Z(_03190_));
 AOI222_X2 _19379_ (.A1(_10778_),
    .A2(_03188_),
    .B1(_03189_),
    .B2(_10794_),
    .C1(_03190_),
    .C2(_10785_),
    .ZN(_03191_));
 NAND2_X1 _19380_ (.A1(_10750_),
    .A2(_03191_),
    .ZN(_03192_));
 MUX2_X1 _19381_ (.A(_01091_),
    .B(_01092_),
    .S(_10628_),
    .Z(_03193_));
 AOI21_X2 _19382_ (.A(_10608_),
    .B1(_03193_),
    .B2(_10616_),
    .ZN(_03194_));
 MUX2_X1 _19383_ (.A(_01087_),
    .B(_01088_),
    .S(_11366_),
    .Z(_03195_));
 AOI21_X2 _19384_ (.A(_11676_),
    .B1(_03195_),
    .B2(_10622_),
    .ZN(_03196_));
 OAI21_X2 _19385_ (.A(_10759_),
    .B1(_03194_),
    .B2(_03196_),
    .ZN(_03197_));
 MUX2_X1 _19386_ (.A(_01085_),
    .B(_01086_),
    .S(_10628_),
    .Z(_03198_));
 INV_X1 _19387_ (.A(_03198_),
    .ZN(_03199_));
 MUX2_X1 _19388_ (.A(_01089_),
    .B(_01090_),
    .S(_10797_),
    .Z(_03200_));
 INV_X1 _19389_ (.A(_03200_),
    .ZN(_03201_));
 AOI221_X2 _19390_ (.A(_10571_),
    .B1(_03196_),
    .B2(_03199_),
    .C1(_03201_),
    .C2(_03194_),
    .ZN(_03202_));
 AOI21_X4 _19391_ (.A(_03192_),
    .B1(_03197_),
    .B2(_03202_),
    .ZN(_03203_));
 OAI21_X2 _19392_ (.A(_11596_),
    .B1(_03185_),
    .B2(_03203_),
    .ZN(_03204_));
 NAND2_X1 _19393_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_10565_),
    .ZN(_03205_));
 INV_X1 _19394_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .ZN(_03206_));
 OAI221_X2 _19395_ (.A(_03204_),
    .B1(_03205_),
    .B2(_10747_),
    .C1(_10673_),
    .C2(_03206_),
    .ZN(_16068_));
 INV_X2 _19396_ (.A(_16068_),
    .ZN(_16072_));
 CLKBUF_X2 _19397_ (.A(_15486_),
    .Z(_03207_));
 INV_X1 _19398_ (.A(_03207_),
    .ZN(_03208_));
 BUF_X2 _19399_ (.A(_15481_),
    .Z(_03209_));
 INV_X1 _19400_ (.A(_15477_),
    .ZN(_03210_));
 AOI21_X1 _19401_ (.A(_15473_),
    .B1(_15469_),
    .B2(_13262_),
    .ZN(_03211_));
 OAI21_X1 _19402_ (.A(_03210_),
    .B1(_03211_),
    .B2(_13260_),
    .ZN(_03212_));
 BUF_X2 _19403_ (.A(_15482_),
    .Z(_03213_));
 AOI21_X1 _19404_ (.A(_03209_),
    .B1(_03212_),
    .B2(_03213_),
    .ZN(_03214_));
 NOR2_X1 _19405_ (.A1(_03208_),
    .A2(_03214_),
    .ZN(_03215_));
 INV_X1 _19406_ (.A(_03213_),
    .ZN(_03216_));
 AOI21_X1 _19407_ (.A(_03216_),
    .B1(_03210_),
    .B2(_13260_),
    .ZN(_03217_));
 NOR3_X2 _19408_ (.A1(_03207_),
    .A2(_03209_),
    .A3(_03217_),
    .ZN(_03218_));
 NOR3_X2 _19409_ (.A1(_13260_),
    .A2(_03216_),
    .A3(_03208_),
    .ZN(_03219_));
 AND3_X2 _19410_ (.A1(_13110_),
    .A2(_13263_),
    .A3(_03219_),
    .ZN(_03220_));
 AOI21_X2 _19411_ (.A(_03209_),
    .B1(_15477_),
    .B2(_03213_),
    .ZN(_03221_));
 NAND3_X1 _19412_ (.A1(_03208_),
    .A2(_03211_),
    .A3(_03221_),
    .ZN(_03222_));
 AOI21_X2 _19413_ (.A(_03222_),
    .B1(_13263_),
    .B2(_13110_),
    .ZN(_03223_));
 NOR4_X4 _19414_ (.A1(_03220_),
    .A2(_03218_),
    .A3(_03215_),
    .A4(_03223_),
    .ZN(\alu_adder_result_ex[29] ));
 OAI21_X1 _19415_ (.A(_15478_),
    .B1(_15473_),
    .B2(_13262_),
    .ZN(_03224_));
 AND3_X1 _19416_ (.A1(_03216_),
    .A2(_03210_),
    .A3(_03224_),
    .ZN(_03225_));
 INV_X1 _19417_ (.A(_15473_),
    .ZN(_03226_));
 OAI21_X2 _19418_ (.A(_03210_),
    .B1(_03226_),
    .B2(_13260_),
    .ZN(_03227_));
 AOI21_X2 _19419_ (.A(_03225_),
    .B1(_03227_),
    .B2(_03213_),
    .ZN(_03228_));
 NAND3_X2 _19420_ (.A1(_13262_),
    .A2(_15478_),
    .A3(_03213_),
    .ZN(_03229_));
 OAI21_X1 _19421_ (.A(_03228_),
    .B1(_03229_),
    .B2(_13275_),
    .ZN(_03230_));
 AOI211_X2 _19422_ (.A(_13272_),
    .B(_03227_),
    .C1(_13274_),
    .C2(_13273_),
    .ZN(_03231_));
 AND2_X1 _19423_ (.A1(_03216_),
    .A2(_03231_),
    .ZN(_03232_));
 NOR3_X1 _19424_ (.A1(_12772_),
    .A2(_03230_),
    .A3(_03232_),
    .ZN(_03233_));
 NAND3_X2 _19425_ (.A1(_12603_),
    .A2(_12605_),
    .A3(_03233_),
    .ZN(_03234_));
 NOR3_X1 _19426_ (.A1(_13267_),
    .A2(_03230_),
    .A3(_03232_),
    .ZN(_03235_));
 AND4_X1 _19427_ (.A1(_12772_),
    .A2(_13267_),
    .A3(_03228_),
    .A4(_03229_),
    .ZN(_03236_));
 NOR2_X1 _19428_ (.A1(_03235_),
    .A2(_03236_),
    .ZN(_03237_));
 NAND3_X2 _19429_ (.A1(_13267_),
    .A2(_03228_),
    .A3(_03229_),
    .ZN(_03238_));
 OAI21_X2 _19430_ (.A(_12602_),
    .B1(_11919_),
    .B2(_11916_),
    .ZN(_03239_));
 OAI211_X4 _19431_ (.A(_03234_),
    .B(_03237_),
    .C1(_03238_),
    .C2(_03239_),
    .ZN(\alu_adder_result_ex[28] ));
 AOI21_X1 _19432_ (.A(_12612_),
    .B1(_11162_),
    .B2(_10498_),
    .ZN(_03240_));
 MUX2_X1 _19433_ (.A(_01100_),
    .B(_01102_),
    .S(_12112_),
    .Z(_03241_));
 NOR2_X1 _19434_ (.A1(_11956_),
    .A2(_03241_),
    .ZN(_03242_));
 MUX2_X1 _19435_ (.A(_01101_),
    .B(_01103_),
    .S(_11978_),
    .Z(_03243_));
 NOR2_X1 _19436_ (.A1(_10697_),
    .A2(_03243_),
    .ZN(_03244_));
 NOR3_X1 _19437_ (.A1(_12029_),
    .A2(_03242_),
    .A3(_03244_),
    .ZN(_03245_));
 INV_X1 _19438_ (.A(_01094_),
    .ZN(_03246_));
 NOR2_X1 _19439_ (.A1(_11952_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .ZN(_03247_));
 AOI21_X1 _19440_ (.A(_03247_),
    .B1(_01095_),
    .B2(_11939_),
    .ZN(_03248_));
 AOI221_X2 _19441_ (.A(_10468_),
    .B1(_03246_),
    .B2(_10964_),
    .C1(_03248_),
    .C2(_12000_),
    .ZN(_03249_));
 NOR3_X2 _19442_ (.A1(_10432_),
    .A2(_03245_),
    .A3(_03249_),
    .ZN(_03250_));
 MUX2_X1 _19443_ (.A(_01104_),
    .B(_01106_),
    .S(_12628_),
    .Z(_03251_));
 MUX2_X1 _19444_ (.A(_01105_),
    .B(_01107_),
    .S(_12628_),
    .Z(_03252_));
 MUX2_X1 _19445_ (.A(_03251_),
    .B(_03252_),
    .S(_12630_),
    .Z(_03253_));
 MUX2_X1 _19446_ (.A(_01096_),
    .B(_01098_),
    .S(_12628_),
    .Z(_03254_));
 MUX2_X1 _19447_ (.A(_01097_),
    .B(_01099_),
    .S(_12704_),
    .Z(_03255_));
 MUX2_X1 _19448_ (.A(_03254_),
    .B(_03255_),
    .S(_12630_),
    .Z(_03256_));
 MUX2_X1 _19449_ (.A(_03253_),
    .B(_03256_),
    .S(_11931_),
    .Z(_03257_));
 NOR2_X1 _19450_ (.A1(_12449_),
    .A2(_03257_),
    .ZN(_03258_));
 NOR3_X2 _19451_ (.A1(_11928_),
    .A2(_03250_),
    .A3(_03258_),
    .ZN(_03259_));
 MUX2_X1 _19452_ (.A(_01116_),
    .B(_01118_),
    .S(_11962_),
    .Z(_03260_));
 MUX2_X1 _19453_ (.A(_01117_),
    .B(_01119_),
    .S(_11938_),
    .Z(_03261_));
 MUX2_X1 _19454_ (.A(_03260_),
    .B(_03261_),
    .S(_12693_),
    .Z(_03262_));
 MUX2_X1 _19455_ (.A(_01108_),
    .B(_01110_),
    .S(net428),
    .Z(_03263_));
 MUX2_X1 _19456_ (.A(_01109_),
    .B(_01111_),
    .S(net427),
    .Z(_03264_));
 MUX2_X1 _19457_ (.A(_03263_),
    .B(_03264_),
    .S(_12693_),
    .Z(_03265_));
 MUX2_X1 _19458_ (.A(_03262_),
    .B(_03265_),
    .S(_11969_),
    .Z(_03266_));
 MUX2_X1 _19459_ (.A(_01120_),
    .B(_01122_),
    .S(net428),
    .Z(_03267_));
 MUX2_X1 _19460_ (.A(_01121_),
    .B(_01123_),
    .S(_12689_),
    .Z(_03268_));
 MUX2_X1 _19461_ (.A(_03267_),
    .B(_03268_),
    .S(_12693_),
    .Z(_03269_));
 MUX2_X1 _19462_ (.A(_01112_),
    .B(_01114_),
    .S(_12689_),
    .Z(_03270_));
 MUX2_X1 _19463_ (.A(_01113_),
    .B(_01115_),
    .S(_12691_),
    .Z(_03271_));
 MUX2_X1 _19464_ (.A(_03270_),
    .B(_03271_),
    .S(_13193_),
    .Z(_03272_));
 MUX2_X1 _19465_ (.A(_03269_),
    .B(_03272_),
    .S(_11969_),
    .Z(_03273_));
 MUX2_X2 _19466_ (.A(_03266_),
    .B(_03273_),
    .S(_12649_),
    .Z(_03274_));
 AOI21_X4 _19467_ (.A(_03259_),
    .B1(_03274_),
    .B2(_11929_),
    .ZN(_03275_));
 OAI21_X1 _19468_ (.A(_11921_),
    .B1(_11994_),
    .B2(_03275_),
    .ZN(_03276_));
 NOR2_X2 _19469_ (.A1(_03240_),
    .A2(_03276_),
    .ZN(_16077_));
 AND3_X1 _19470_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(_10564_),
    .A3(_10870_),
    .ZN(_03277_));
 MUX2_X1 _19471_ (.A(_01100_),
    .B(_01102_),
    .S(_11454_),
    .Z(_03278_));
 NOR2_X1 _19472_ (.A1(_10628_),
    .A2(_03278_),
    .ZN(_03279_));
 MUX2_X1 _19473_ (.A(_01101_),
    .B(_01103_),
    .S(_11363_),
    .Z(_03280_));
 NOR2_X1 _19474_ (.A1(_10580_),
    .A2(_03280_),
    .ZN(_03281_));
 NOR3_X1 _19475_ (.A1(_10828_),
    .A2(_03279_),
    .A3(_03281_),
    .ZN(_03282_));
 NOR2_X1 _19476_ (.A1(_10613_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .ZN(_03283_));
 AOI21_X1 _19477_ (.A(_03283_),
    .B1(_01095_),
    .B2(_10587_),
    .ZN(_03284_));
 AOI221_X2 _19478_ (.A(_10765_),
    .B1(_03246_),
    .B2(_10822_),
    .C1(_03284_),
    .C2(_10796_),
    .ZN(_03285_));
 NOR3_X2 _19479_ (.A1(_11676_),
    .A2(_03282_),
    .A3(_03285_),
    .ZN(_03286_));
 MUX2_X1 _19480_ (.A(_01104_),
    .B(_01106_),
    .S(_11642_),
    .Z(_03287_));
 MUX2_X1 _19481_ (.A(_01105_),
    .B(_01107_),
    .S(_11642_),
    .Z(_03288_));
 MUX2_X1 _19482_ (.A(_03287_),
    .B(_03288_),
    .S(_10862_),
    .Z(_03289_));
 MUX2_X1 _19483_ (.A(_01096_),
    .B(_01098_),
    .S(_11642_),
    .Z(_03290_));
 MUX2_X1 _19484_ (.A(_01097_),
    .B(_01099_),
    .S(_11642_),
    .Z(_03291_));
 MUX2_X1 _19485_ (.A(_03290_),
    .B(_03291_),
    .S(_10862_),
    .Z(_03292_));
 MUX2_X1 _19486_ (.A(_03289_),
    .B(_03292_),
    .S(_11357_),
    .Z(_03293_));
 NOR2_X1 _19487_ (.A1(_10608_),
    .A2(_03293_),
    .ZN(_03294_));
 NOR3_X2 _19488_ (.A1(_10749_),
    .A2(_03286_),
    .A3(_03294_),
    .ZN(_03295_));
 MUX2_X1 _19489_ (.A(_01116_),
    .B(_01118_),
    .S(_11771_),
    .Z(_03296_));
 MUX2_X1 _19490_ (.A(_01117_),
    .B(_01119_),
    .S(_11771_),
    .Z(_03297_));
 MUX2_X1 _19491_ (.A(_03296_),
    .B(_03297_),
    .S(_11534_),
    .Z(_03298_));
 MUX2_X1 _19492_ (.A(_01108_),
    .B(_01110_),
    .S(_11771_),
    .Z(_03299_));
 MUX2_X1 _19493_ (.A(_01109_),
    .B(_01111_),
    .S(_11771_),
    .Z(_03300_));
 MUX2_X1 _19494_ (.A(_03299_),
    .B(_03300_),
    .S(_11534_),
    .Z(_03301_));
 MUX2_X1 _19495_ (.A(_03298_),
    .B(_03301_),
    .S(_10569_),
    .Z(_03302_));
 MUX2_X1 _19496_ (.A(_01120_),
    .B(_01122_),
    .S(_11771_),
    .Z(_03303_));
 MUX2_X1 _19497_ (.A(_01121_),
    .B(_01123_),
    .S(_12317_),
    .Z(_03304_));
 MUX2_X1 _19498_ (.A(_03303_),
    .B(_03304_),
    .S(_10627_),
    .Z(_03305_));
 MUX2_X1 _19499_ (.A(_01112_),
    .B(_01114_),
    .S(_11771_),
    .Z(_03306_));
 MUX2_X1 _19500_ (.A(_01113_),
    .B(_01115_),
    .S(_12317_),
    .Z(_03307_));
 MUX2_X1 _19501_ (.A(_03306_),
    .B(_03307_),
    .S(_10627_),
    .Z(_03308_));
 MUX2_X1 _19502_ (.A(_03305_),
    .B(_03308_),
    .S(_10828_),
    .Z(_03309_));
 MUX2_X2 _19503_ (.A(_03302_),
    .B(_03309_),
    .S(_10752_),
    .Z(_03310_));
 AOI21_X4 _19504_ (.A(_03295_),
    .B1(_03310_),
    .B2(_10750_),
    .ZN(_03311_));
 AOI221_X2 _19505_ (.A(_03277_),
    .B1(_03311_),
    .B2(_11596_),
    .C1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .C2(_10397_),
    .ZN(_03312_));
 BUF_X4 _19506_ (.A(_03312_),
    .Z(_16080_));
 AOI221_X2 _19507_ (.A(_10403_),
    .B1(_10928_),
    .B2(_11320_),
    .C1(_10930_),
    .C2(_10509_),
    .ZN(_03313_));
 MUX2_X1 _19508_ (.A(_01147_),
    .B(_01149_),
    .S(_10452_),
    .Z(_03314_));
 MUX2_X1 _19509_ (.A(_01148_),
    .B(_01150_),
    .S(_10452_),
    .Z(_03315_));
 MUX2_X1 _19510_ (.A(_03314_),
    .B(_03315_),
    .S(_10941_),
    .Z(_03316_));
 MUX2_X1 _19511_ (.A(_01139_),
    .B(_01141_),
    .S(_10452_),
    .Z(_03317_));
 MUX2_X1 _19512_ (.A(_01140_),
    .B(_01142_),
    .S(_10452_),
    .Z(_03318_));
 MUX2_X1 _19513_ (.A(_03317_),
    .B(_03318_),
    .S(_10941_),
    .Z(_03319_));
 MUX2_X1 _19514_ (.A(_03316_),
    .B(_03319_),
    .S(_10421_),
    .Z(_03320_));
 NAND3_X2 _19515_ (.A1(_10435_),
    .A2(_10709_),
    .A3(_03320_),
    .ZN(_03321_));
 MUX2_X1 _19516_ (.A(_01144_),
    .B(_01146_),
    .S(_10437_),
    .Z(_03322_));
 NOR2_X1 _19517_ (.A1(_10695_),
    .A2(_03322_),
    .ZN(_03323_));
 MUX2_X1 _19518_ (.A(_01143_),
    .B(_01145_),
    .S(_10456_),
    .Z(_03324_));
 NOR2_X1 _19519_ (.A1(_10442_),
    .A2(_03324_),
    .ZN(_03325_));
 NOR2_X1 _19520_ (.A1(_10452_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .ZN(_03326_));
 AND2_X1 _19521_ (.A1(_10437_),
    .A2(_01126_),
    .ZN(_03327_));
 NOR3_X1 _19522_ (.A1(_10695_),
    .A2(_03326_),
    .A3(_03327_),
    .ZN(_03328_));
 NOR3_X1 _19523_ (.A1(_10879_),
    .A2(_10337_),
    .A3(_01125_),
    .ZN(_03329_));
 OAI33_X1 _19524_ (.A1(_11099_),
    .A2(_03323_),
    .A3(_03325_),
    .B1(_03328_),
    .B2(_03329_),
    .B3(_10998_),
    .ZN(_03330_));
 MUX2_X1 _19525_ (.A(_01152_),
    .B(_01154_),
    .S(net334),
    .Z(_03331_));
 NOR2_X1 _19526_ (.A1(_10695_),
    .A2(_03331_),
    .ZN(_03332_));
 MUX2_X1 _19527_ (.A(_01151_),
    .B(_01153_),
    .S(net334),
    .Z(_03333_));
 NOR2_X1 _19528_ (.A1(_10442_),
    .A2(_03333_),
    .ZN(_03334_));
 MUX2_X1 _19529_ (.A(_01127_),
    .B(_01129_),
    .S(_10408_),
    .Z(_03335_));
 NOR2_X1 _19530_ (.A1(_10442_),
    .A2(_03335_),
    .ZN(_03336_));
 MUX2_X1 _19531_ (.A(_01128_),
    .B(_01130_),
    .S(_10408_),
    .Z(_03337_));
 NOR2_X1 _19532_ (.A1(_10694_),
    .A2(_03337_),
    .ZN(_03338_));
 NAND2_X1 _19533_ (.A1(_10420_),
    .A2(_10472_),
    .ZN(_03339_));
 OAI33_X1 _19534_ (.A1(_11042_),
    .A2(_03332_),
    .A3(_03334_),
    .B1(_03336_),
    .B2(_03338_),
    .B3(_03339_),
    .ZN(_03340_));
 MUX2_X1 _19535_ (.A(_01134_),
    .B(_01138_),
    .S(_10978_),
    .Z(_03341_));
 NOR2_X1 _19536_ (.A1(_10977_),
    .A2(_03341_),
    .ZN(_03342_));
 MUX2_X1 _19537_ (.A(_01132_),
    .B(_01136_),
    .S(_10434_),
    .Z(_03343_));
 NOR3_X1 _19538_ (.A1(_11186_),
    .A2(net397),
    .A3(_03343_),
    .ZN(_03344_));
 MUX2_X1 _19539_ (.A(_01131_),
    .B(_01135_),
    .S(_10684_),
    .Z(_03345_));
 NOR2_X1 _19540_ (.A1(_10980_),
    .A2(_03345_),
    .ZN(_03346_));
 NOR3_X1 _19541_ (.A1(_03342_),
    .A2(_03344_),
    .A3(_03346_),
    .ZN(_03347_));
 MUX2_X1 _19542_ (.A(_01133_),
    .B(_01137_),
    .S(_10684_),
    .Z(_03348_));
 NOR3_X1 _19543_ (.A1(_10941_),
    .A2(_10337_),
    .A3(_03348_),
    .ZN(_03349_));
 NOR2_X1 _19544_ (.A1(_10962_),
    .A2(_03349_),
    .ZN(_03350_));
 AOI221_X2 _19545_ (.A(_03330_),
    .B1(_03340_),
    .B2(_10432_),
    .C1(_03347_),
    .C2(_03350_),
    .ZN(_03351_));
 AOI21_X1 _19546_ (.A(_10317_),
    .B1(_03321_),
    .B2(_03351_),
    .ZN(_03352_));
 OR2_X2 _19547_ (.A1(_10361_),
    .A2(_03352_),
    .ZN(_03353_));
 NOR2_X2 _19548_ (.A1(_03313_),
    .A2(_03353_),
    .ZN(_15495_));
 NAND2_X1 _19549_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(_10361_),
    .ZN(_03354_));
 INV_X1 _19550_ (.A(_01125_),
    .ZN(_03355_));
 NOR2_X1 _19551_ (.A1(_10857_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .ZN(_03356_));
 AOI21_X1 _19552_ (.A(_03356_),
    .B1(_01126_),
    .B2(_11567_),
    .ZN(_03357_));
 AOI221_X2 _19553_ (.A(_10764_),
    .B1(_03355_),
    .B2(_10821_),
    .C1(_03357_),
    .C2(_10861_),
    .ZN(_03358_));
 MUX2_X1 _19554_ (.A(_01131_),
    .B(_01133_),
    .S(_10598_),
    .Z(_03359_));
 NAND3_X1 _19555_ (.A1(_10579_),
    .A2(_10765_),
    .A3(_03359_),
    .ZN(_03360_));
 MUX2_X1 _19556_ (.A(_01132_),
    .B(_01134_),
    .S(_10857_),
    .Z(_03361_));
 NAND3_X1 _19557_ (.A1(_10786_),
    .A2(_10764_),
    .A3(_03361_),
    .ZN(_03362_));
 NAND4_X2 _19558_ (.A1(_10607_),
    .A2(_10573_),
    .A3(_03360_),
    .A4(_03362_),
    .ZN(_03363_));
 MUX2_X1 _19559_ (.A(_01135_),
    .B(_01137_),
    .S(_10856_),
    .Z(_03364_));
 MUX2_X1 _19560_ (.A(_01136_),
    .B(_01138_),
    .S(_10856_),
    .Z(_03365_));
 MUX2_X1 _19561_ (.A(_03364_),
    .B(_03365_),
    .S(_10592_),
    .Z(_03366_));
 MUX2_X1 _19562_ (.A(_01127_),
    .B(_01129_),
    .S(_10856_),
    .Z(_03367_));
 MUX2_X1 _19563_ (.A(_01128_),
    .B(_01130_),
    .S(_10856_),
    .Z(_03368_));
 MUX2_X1 _19564_ (.A(_03367_),
    .B(_03368_),
    .S(_10592_),
    .Z(_03369_));
 MUX2_X1 _19565_ (.A(_03366_),
    .B(_03369_),
    .S(_10567_),
    .Z(_03370_));
 OAI22_X4 _19566_ (.A1(_03358_),
    .A2(_03363_),
    .B1(_03370_),
    .B2(_10855_),
    .ZN(_03371_));
 MUX2_X1 _19567_ (.A(_01144_),
    .B(_01146_),
    .S(_10584_),
    .Z(_03372_));
 MUX2_X1 _19568_ (.A(_01143_),
    .B(_01145_),
    .S(_10584_),
    .Z(_03373_));
 MUX2_X1 _19569_ (.A(_03372_),
    .B(_03373_),
    .S(_10578_),
    .Z(_03374_));
 MUX2_X1 _19570_ (.A(_01141_),
    .B(_01142_),
    .S(_10592_),
    .Z(_03375_));
 AOI22_X1 _19571_ (.A1(_10778_),
    .A2(_03374_),
    .B1(_03375_),
    .B2(_10793_),
    .ZN(_03376_));
 MUX2_X1 _19572_ (.A(_01139_),
    .B(_01140_),
    .S(_10625_),
    .Z(_03377_));
 AOI21_X1 _19573_ (.A(_10573_),
    .B1(_10784_),
    .B2(_03377_),
    .ZN(_03378_));
 MUX2_X1 _19574_ (.A(_01151_),
    .B(_01153_),
    .S(_10584_),
    .Z(_03379_));
 MUX2_X1 _19575_ (.A(_01152_),
    .B(_01154_),
    .S(_10584_),
    .Z(_03380_));
 MUX2_X1 _19576_ (.A(_03379_),
    .B(_03380_),
    .S(_10592_),
    .Z(_03381_));
 MUX2_X1 _19577_ (.A(_01147_),
    .B(_01149_),
    .S(_10856_),
    .Z(_03382_));
 MUX2_X1 _19578_ (.A(_01148_),
    .B(_01150_),
    .S(_10856_),
    .Z(_03383_));
 MUX2_X1 _19579_ (.A(_03382_),
    .B(_03383_),
    .S(_10592_),
    .Z(_03384_));
 AOI22_X1 _19580_ (.A1(_10651_),
    .A2(_03381_),
    .B1(_03384_),
    .B2(_10643_),
    .ZN(_03385_));
 AND3_X2 _19581_ (.A1(_03376_),
    .A2(_03378_),
    .A3(_03385_),
    .ZN(_03386_));
 OAI221_X2 _19582_ (.A(_10563_),
    .B1(_03371_),
    .B2(_03386_),
    .C1(_10681_),
    .C2(_10361_),
    .ZN(_03387_));
 NAND4_X2 _19583_ (.A1(\cs_registers_i.pc_id_i[31] ),
    .A2(_10326_),
    .A3(_10563_),
    .A4(_10672_),
    .ZN(_03388_));
 NAND3_X4 _19584_ (.A1(_03354_),
    .A2(_03387_),
    .A3(_03388_),
    .ZN(_15496_));
 INV_X2 _19585_ (.A(_15496_),
    .ZN(_15492_));
 AND2_X1 _19586_ (.A1(_15490_),
    .A2(_03219_),
    .ZN(_03389_));
 INV_X1 _19587_ (.A(_15485_),
    .ZN(_03390_));
 OAI21_X2 _19588_ (.A(_03390_),
    .B1(_03221_),
    .B2(_03208_),
    .ZN(_03391_));
 AOI221_X2 _19589_ (.A(_15489_),
    .B1(_13266_),
    .B2(_03389_),
    .C1(_03391_),
    .C2(_15490_),
    .ZN(_03392_));
 NOR2_X1 _19590_ (.A1(_11632_),
    .A2(_03352_),
    .ZN(_03393_));
 NAND3_X1 _19591_ (.A1(_10503_),
    .A2(_10389_),
    .A3(_10928_),
    .ZN(_03394_));
 OAI221_X2 _19592_ (.A(_10317_),
    .B1(_10926_),
    .B2(_03394_),
    .C1(_10387_),
    .C2(_10510_),
    .ZN(_03395_));
 AOI21_X4 _19593_ (.A(_15496_),
    .B1(_03393_),
    .B2(_03395_),
    .ZN(_03396_));
 NOR3_X4 _19594_ (.A1(_03313_),
    .A2(_03353_),
    .A3(_15492_),
    .ZN(_03397_));
 OAI21_X4 _19595_ (.A(_11514_),
    .B1(_03396_),
    .B2(_03397_),
    .ZN(_03398_));
 OR4_X4 _19596_ (.A1(_11401_),
    .A2(_11863_),
    .A3(_03396_),
    .A4(_03397_),
    .ZN(_03399_));
 NAND2_X2 _19597_ (.A1(_03321_),
    .A2(_03351_),
    .ZN(_03400_));
 BUF_X2 _19598_ (.A(_00179_),
    .Z(_03401_));
 BUF_X4 _19599_ (.A(_00178_),
    .Z(_03402_));
 BUF_X4 _19600_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Z(_03403_));
 BUF_X4 _19601_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Z(_03404_));
 NOR2_X4 _19602_ (.A1(_03403_),
    .A2(_03404_),
    .ZN(_03405_));
 NAND3_X4 _19603_ (.A1(_03401_),
    .A2(_03402_),
    .A3(_03405_),
    .ZN(_03406_));
 INV_X4 _19604_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .ZN(_03407_));
 CLKBUF_X3 _19605_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .Z(_03408_));
 OAI221_X2 _19606_ (.A(_03406_),
    .B1(_03405_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .C1(_03407_),
    .C2(_03408_),
    .ZN(_03409_));
 NOR3_X1 _19607_ (.A1(_03402_),
    .A2(_03371_),
    .A3(_03386_),
    .ZN(_03410_));
 OAI22_X2 _19608_ (.A1(_03400_),
    .A2(_03406_),
    .B1(_03409_),
    .B2(_03410_),
    .ZN(_03411_));
 CLKBUF_X3 _19609_ (.A(_01155_),
    .Z(_03412_));
 NOR2_X1 _19610_ (.A1(_03412_),
    .A2(_03405_),
    .ZN(_03413_));
 XNOR2_X1 _19611_ (.A(_03411_),
    .B(_03413_),
    .ZN(_03414_));
 OR2_X2 _19612_ (.A1(_11405_),
    .A2(_03414_),
    .ZN(_03415_));
 NAND3_X4 _19613_ (.A1(_03398_),
    .A2(_03399_),
    .A3(_03415_),
    .ZN(_03416_));
 XNOR2_X2 _19614_ (.A(_03392_),
    .B(_03416_),
    .ZN(_03417_));
 INV_X4 _19615_ (.A(_03417_),
    .ZN(\alu_adder_result_ex[31] ));
 INV_X2 _19616_ (.A(_15490_),
    .ZN(_03418_));
 NOR3_X1 _19617_ (.A1(_03418_),
    .A2(_03209_),
    .A3(_15485_),
    .ZN(_03419_));
 NAND2_X1 _19618_ (.A1(_13099_),
    .A2(_13107_),
    .ZN(_03420_));
 OAI211_X2 _19619_ (.A(_03231_),
    .B(_03419_),
    .C1(_12610_),
    .C2(_03420_),
    .ZN(_03421_));
 AOI21_X1 _19620_ (.A(_03216_),
    .B1(_03210_),
    .B2(_03224_),
    .ZN(_03422_));
 OAI21_X1 _19621_ (.A(_03207_),
    .B1(_03209_),
    .B2(_03422_),
    .ZN(_03423_));
 AOI21_X1 _19622_ (.A(_03418_),
    .B1(_03390_),
    .B2(_03423_),
    .ZN(_03424_));
 AOI21_X1 _19623_ (.A(_15485_),
    .B1(_03209_),
    .B2(_03207_),
    .ZN(_03425_));
 AND2_X1 _19624_ (.A1(_03418_),
    .A2(_03425_),
    .ZN(_03426_));
 NAND3_X1 _19625_ (.A1(_03207_),
    .A2(_03418_),
    .A3(_03422_),
    .ZN(_03427_));
 INV_X1 _19626_ (.A(_03231_),
    .ZN(_03428_));
 AOI21_X1 _19627_ (.A(_03428_),
    .B1(_13267_),
    .B2(_13119_),
    .ZN(_03429_));
 OAI221_X2 _19628_ (.A(_03421_),
    .B1(_03424_),
    .B2(_03426_),
    .C1(_03427_),
    .C2(_03429_),
    .ZN(_03430_));
 BUF_X8 _19629_ (.A(_03430_),
    .Z(\alu_adder_result_ex[30] ));
 BUF_X4 _19630_ (.A(_03403_),
    .Z(_03431_));
 INV_X2 _19631_ (.A(_03431_),
    .ZN(_03432_));
 OR4_X2 _19632_ (.A1(_10894_),
    .A2(_10910_),
    .A3(_10918_),
    .A4(_11417_),
    .ZN(_03433_));
 BUF_X8 _19633_ (.A(_03433_),
    .Z(_03434_));
 INV_X2 _19634_ (.A(_11419_),
    .ZN(_03435_));
 INV_X4 _19635_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_03436_));
 NOR4_X4 _19636_ (.A1(_03436_),
    .A2(_11421_),
    .A3(_11422_),
    .A4(_11424_),
    .ZN(_03437_));
 NAND3_X4 _19637_ (.A1(_10304_),
    .A2(_03435_),
    .A3(_03437_),
    .ZN(_03438_));
 NOR2_X4 _19638_ (.A1(_03434_),
    .A2(_03438_),
    .ZN(_03439_));
 NOR2_X4 _19639_ (.A1(_12103_),
    .A2(_11407_),
    .ZN(_03440_));
 NAND2_X4 _19640_ (.A1(_03439_),
    .A2(_03440_),
    .ZN(_03441_));
 BUF_X2 _19641_ (.A(_01158_),
    .Z(_03442_));
 AND2_X1 _19642_ (.A1(_03442_),
    .A2(_15546_),
    .ZN(_03443_));
 CLKBUF_X2 _19643_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .Z(_03444_));
 CLKBUF_X3 _19644_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Z(_03445_));
 NOR2_X1 _19645_ (.A1(_03444_),
    .A2(_03445_),
    .ZN(_03446_));
 NAND2_X1 _19646_ (.A1(_03443_),
    .A2(_03446_),
    .ZN(_03447_));
 OR3_X1 _19647_ (.A1(_03432_),
    .A2(_03441_),
    .A3(_03447_),
    .ZN(_03448_));
 BUF_X4 _19648_ (.A(_11401_),
    .Z(_03449_));
 NAND2_X4 _19649_ (.A1(net300),
    .A2(_03449_),
    .ZN(_03450_));
 NOR2_X4 _19650_ (.A1(_11428_),
    .A2(_03450_),
    .ZN(_03451_));
 INV_X1 _19651_ (.A(_03404_),
    .ZN(_03452_));
 OAI21_X1 _19652_ (.A(_03448_),
    .B1(_03451_),
    .B2(_03452_),
    .ZN(_00002_));
 CLKBUF_X3 _19653_ (.A(data_rvalid_i),
    .Z(_03453_));
 NOR2_X4 _19654_ (.A1(_10324_),
    .A2(net302),
    .ZN(_03454_));
 AND2_X2 _19655_ (.A1(_10320_),
    .A2(_03454_),
    .ZN(_03455_));
 NAND2_X2 _19656_ (.A1(_03453_),
    .A2(_03455_),
    .ZN(_03456_));
 NOR2_X2 _19657_ (.A1(net36),
    .A2(\load_store_unit_i.lsu_err_q ),
    .ZN(_03457_));
 NOR3_X2 _19658_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_03456_),
    .A3(_03457_),
    .ZN(\id_stage_i.controller_i.load_err_d ));
 NOR3_X2 _19659_ (.A1(_01160_),
    .A2(_03456_),
    .A3(_03457_),
    .ZN(\id_stage_i.controller_i.store_err_d ));
 INV_X4 _19660_ (.A(_11421_),
    .ZN(_03458_));
 NOR3_X4 _19661_ (.A1(_03458_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A3(_11424_),
    .ZN(_03459_));
 AND2_X1 _19662_ (.A1(_03436_),
    .A2(_03459_),
    .ZN(_03460_));
 BUF_X4 _19663_ (.A(_03460_),
    .Z(_03461_));
 BUF_X1 _19664_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .Z(_03462_));
 BUF_X1 _19665_ (.A(\cs_registers_i.priv_lvl_q[1] ),
    .Z(_03463_));
 AND2_X1 _19666_ (.A1(_03462_),
    .A2(_03463_),
    .ZN(_03464_));
 BUF_X4 _19667_ (.A(_10557_),
    .Z(_03465_));
 NOR2_X2 _19668_ (.A1(_03465_),
    .A2(_10876_),
    .ZN(_03466_));
 NAND3_X4 _19669_ (.A1(_10304_),
    .A2(_10522_),
    .A3(_10670_),
    .ZN(_03467_));
 NOR3_X4 _19670_ (.A1(_10891_),
    .A2(_10886_),
    .A3(_03467_),
    .ZN(_03468_));
 AND2_X2 _19671_ (.A1(_03466_),
    .A2(_03468_),
    .ZN(_03469_));
 OR3_X2 _19672_ (.A1(_10878_),
    .A2(_10880_),
    .A3(_10881_),
    .ZN(_03470_));
 OR2_X2 _19673_ (.A1(_03465_),
    .A2(_10876_),
    .ZN(_03471_));
 NOR4_X4 _19674_ (.A1(_01161_),
    .A2(_10742_),
    .A3(_03470_),
    .A4(_03471_),
    .ZN(_03472_));
 AOI21_X1 _19675_ (.A(_03469_),
    .B1(_03472_),
    .B2(\cs_registers_i.csr_mstatus_tw_o ),
    .ZN(_03473_));
 NOR2_X1 _19676_ (.A1(_03464_),
    .A2(_03473_),
    .ZN(_03474_));
 NOR2_X2 _19677_ (.A1(_10887_),
    .A2(_10889_),
    .ZN(_03475_));
 AND3_X2 _19678_ (.A1(_10661_),
    .A2(_03475_),
    .A3(_03468_),
    .ZN(_03476_));
 CLKBUF_X3 _19679_ (.A(\cs_registers_i.debug_mode_i ),
    .Z(_03477_));
 INV_X2 _19680_ (.A(_03477_),
    .ZN(_03478_));
 AOI21_X2 _19681_ (.A(_03474_),
    .B1(_03476_),
    .B2(_03478_),
    .ZN(_03479_));
 INV_X1 _19682_ (.A(_03479_),
    .ZN(_03480_));
 NAND2_X1 _19683_ (.A1(_15502_),
    .A2(_15505_),
    .ZN(_03481_));
 INV_X1 _19684_ (.A(_15502_),
    .ZN(_03482_));
 NOR2_X1 _19685_ (.A1(_03482_),
    .A2(_15504_),
    .ZN(_03483_));
 OAI21_X2 _19686_ (.A(_03481_),
    .B1(_03483_),
    .B2(_15501_),
    .ZN(_03484_));
 NOR3_X4 _19687_ (.A1(_15920_),
    .A2(_11321_),
    .A3(_11352_),
    .ZN(_03485_));
 NAND2_X1 _19688_ (.A1(_10921_),
    .A2(_11427_),
    .ZN(_03486_));
 NOR2_X1 _19689_ (.A1(_15527_),
    .A2(_03486_),
    .ZN(_03487_));
 NAND2_X1 _19690_ (.A1(_03485_),
    .A2(_03487_),
    .ZN(_03488_));
 NOR2_X2 _19691_ (.A1(_10744_),
    .A2(_03434_),
    .ZN(_03489_));
 OAI33_X1 _19692_ (.A1(_10885_),
    .A2(_10923_),
    .A3(_11074_),
    .B1(_11241_),
    .B2(_11279_),
    .B3(_10974_),
    .ZN(_03490_));
 BUF_X4 _19693_ (.A(_03490_),
    .Z(_03491_));
 AND4_X1 _19694_ (.A1(_03489_),
    .A2(_15916_),
    .A3(_15929_),
    .A4(_03491_),
    .ZN(_03492_));
 NOR2_X4 _19695_ (.A1(_03465_),
    .A2(_10678_),
    .ZN(_03493_));
 NAND2_X1 _19696_ (.A1(_03493_),
    .A2(_11418_),
    .ZN(_03494_));
 BUF_X4 _19697_ (.A(_03494_),
    .Z(_03495_));
 NOR2_X2 _19698_ (.A1(_11065_),
    .A2(_03495_),
    .ZN(_03496_));
 NOR2_X1 _19699_ (.A1(_15884_),
    .A2(_15896_),
    .ZN(_03497_));
 NAND4_X4 _19700_ (.A1(_15876_),
    .A2(_03492_),
    .A3(_03496_),
    .A4(_03497_),
    .ZN(_03498_));
 BUF_X4 _19701_ (.A(_03495_),
    .Z(_03499_));
 INV_X4 _19702_ (.A(_15515_),
    .ZN(_03500_));
 BUF_X4 _19703_ (.A(_15512_),
    .Z(_03501_));
 INV_X4 _19704_ (.A(_03501_),
    .ZN(_03502_));
 CLKBUF_X3 _19705_ (.A(_15520_),
    .Z(_03503_));
 INV_X2 _19706_ (.A(_03503_),
    .ZN(_03504_));
 NAND3_X4 _19707_ (.A1(_03500_),
    .A2(_03502_),
    .A3(_03504_),
    .ZN(_03505_));
 BUF_X4 _19708_ (.A(_15518_),
    .Z(_03506_));
 OAI221_X2 _19709_ (.A(_03478_),
    .B1(_11071_),
    .B2(_03499_),
    .C1(_03505_),
    .C2(_03506_),
    .ZN(_03507_));
 OAI211_X4 _19710_ (.A(_03484_),
    .B(_03488_),
    .C1(_03498_),
    .C2(_03507_),
    .ZN(_03508_));
 AOI21_X2 _19711_ (.A(_03434_),
    .B1(_03508_),
    .B2(_03493_),
    .ZN(_03509_));
 INV_X2 _19712_ (.A(_15518_),
    .ZN(_03510_));
 NOR3_X1 _19713_ (.A1(_11066_),
    .A2(_03501_),
    .A3(_03503_),
    .ZN(_03511_));
 NAND2_X1 _19714_ (.A1(_03510_),
    .A2(_03511_),
    .ZN(_03512_));
 NAND2_X2 _19715_ (.A1(_15888_),
    .A2(_15896_),
    .ZN(_03513_));
 NOR2_X4 _19716_ (.A1(_15876_),
    .A2(_03513_),
    .ZN(_03514_));
 NAND2_X2 _19717_ (.A1(_15920_),
    .A2(_03491_),
    .ZN(_03515_));
 NOR3_X1 _19718_ (.A1(_03495_),
    .A2(_15929_),
    .A3(_03515_),
    .ZN(_03516_));
 AND4_X1 _19719_ (.A1(_03512_),
    .A2(_03496_),
    .A3(_03514_),
    .A4(_03516_),
    .ZN(_03517_));
 BUF_X4 _19720_ (.A(_03489_),
    .Z(_03518_));
 AND4_X4 _19721_ (.A1(_11033_),
    .A2(_11041_),
    .A3(_11049_),
    .A4(_11056_),
    .ZN(_03519_));
 INV_X1 _19722_ (.A(_00138_),
    .ZN(_03520_));
 MUX2_X1 _19723_ (.A(_03520_),
    .B(_11928_),
    .S(_10386_),
    .Z(_03521_));
 AOI22_X2 _19724_ (.A1(_10976_),
    .A2(_03519_),
    .B1(_03521_),
    .B2(_11020_),
    .ZN(_03522_));
 OAI211_X2 _19725_ (.A(_10903_),
    .B(_10386_),
    .C1(_10387_),
    .C2(_10392_),
    .ZN(_03523_));
 NAND3_X2 _19726_ (.A1(_03522_),
    .A2(_03523_),
    .A3(_15880_),
    .ZN(_03524_));
 OAI21_X1 _19727_ (.A(_03518_),
    .B1(_03513_),
    .B2(_03524_),
    .ZN(_03525_));
 AND2_X1 _19728_ (.A1(_03525_),
    .A2(_03516_),
    .ZN(_03526_));
 NOR3_X2 _19729_ (.A1(_11066_),
    .A2(_03506_),
    .A3(_03503_),
    .ZN(_03527_));
 NAND2_X1 _19730_ (.A1(_03499_),
    .A2(_03527_),
    .ZN(_03528_));
 NAND2_X1 _19731_ (.A1(_03512_),
    .A2(_03528_),
    .ZN(_03529_));
 BUF_X4 _19732_ (.A(_11071_),
    .Z(_03530_));
 AOI21_X2 _19733_ (.A(_03529_),
    .B1(_03527_),
    .B2(_03530_),
    .ZN(_03531_));
 AOI21_X4 _19734_ (.A(_03517_),
    .B1(_03526_),
    .B2(_03531_),
    .ZN(_03532_));
 NOR2_X2 _19735_ (.A1(_15929_),
    .A2(_03515_),
    .ZN(_03533_));
 OAI21_X2 _19736_ (.A(_11159_),
    .B1(_11160_),
    .B2(_11162_),
    .ZN(_03534_));
 NOR3_X1 _19737_ (.A1(_03495_),
    .A2(_03534_),
    .A3(_15896_),
    .ZN(_03535_));
 NAND2_X1 _19738_ (.A1(_03533_),
    .A2(_03535_),
    .ZN(_03536_));
 NOR3_X4 _19739_ (.A1(_11061_),
    .A2(_11063_),
    .A3(_11116_),
    .ZN(_03537_));
 OAI22_X1 _19740_ (.A1(_11066_),
    .A2(_03503_),
    .B1(_03495_),
    .B2(_03537_),
    .ZN(_03538_));
 OAI21_X2 _19741_ (.A(_11025_),
    .B1(_10975_),
    .B2(_10934_),
    .ZN(_03539_));
 BUF_X4 _19742_ (.A(_03539_),
    .Z(_03540_));
 AOI21_X1 _19743_ (.A(_03538_),
    .B1(_03518_),
    .B2(_03540_),
    .ZN(_03541_));
 NOR2_X1 _19744_ (.A1(_10919_),
    .A2(_15876_),
    .ZN(_03542_));
 NAND2_X1 _19745_ (.A1(_15869_),
    .A2(_03542_),
    .ZN(_03543_));
 OAI33_X1 _19746_ (.A1(_11066_),
    .A2(_03501_),
    .A3(_03503_),
    .B1(_10934_),
    .B2(_10975_),
    .B3(_15864_),
    .ZN(_03544_));
 AOI221_X1 _19747_ (.A(_03543_),
    .B1(_03511_),
    .B2(_11071_),
    .C1(_03510_),
    .C2(_03544_),
    .ZN(_03545_));
 NAND2_X1 _19748_ (.A1(_03489_),
    .A2(_03505_),
    .ZN(_03546_));
 OAI21_X1 _19749_ (.A(_03510_),
    .B1(_11071_),
    .B2(_03546_),
    .ZN(_03547_));
 NOR4_X1 _19750_ (.A1(_10934_),
    .A2(_10975_),
    .A3(_11065_),
    .A4(_03505_),
    .ZN(_03548_));
 OAI21_X1 _19751_ (.A(_15880_),
    .B1(_11065_),
    .B2(_15860_),
    .ZN(_03549_));
 OAI21_X1 _19752_ (.A(_03518_),
    .B1(_03548_),
    .B2(_03549_),
    .ZN(_03550_));
 AOI211_X4 _19753_ (.A(_03541_),
    .B(_03545_),
    .C1(_03547_),
    .C2(_03550_),
    .ZN(_03551_));
 OAI211_X2 _19754_ (.A(_03493_),
    .B(_03532_),
    .C1(_03536_),
    .C2(_03551_),
    .ZN(_03552_));
 NOR3_X4 _19755_ (.A1(_03495_),
    .A2(_15925_),
    .A3(_03515_),
    .ZN(_03553_));
 NOR3_X2 _19756_ (.A1(_10919_),
    .A2(_15884_),
    .A3(_15896_),
    .ZN(_03554_));
 NOR2_X1 _19757_ (.A1(_15518_),
    .A2(_03505_),
    .ZN(_03555_));
 NOR2_X1 _19758_ (.A1(_15880_),
    .A2(_03555_),
    .ZN(_03556_));
 NAND3_X1 _19759_ (.A1(_15869_),
    .A2(_03554_),
    .A3(_03556_),
    .ZN(_03557_));
 NOR3_X1 _19760_ (.A1(_10920_),
    .A2(_03530_),
    .A3(_03557_),
    .ZN(_03558_));
 NOR4_X1 _19761_ (.A1(_11061_),
    .A2(_11063_),
    .A3(_15876_),
    .A4(_15892_),
    .ZN(_03559_));
 OAI21_X1 _19762_ (.A(_11066_),
    .B1(_03499_),
    .B2(_03559_),
    .ZN(_03560_));
 AOI21_X1 _19763_ (.A(_03560_),
    .B1(_03518_),
    .B2(_03540_),
    .ZN(_03561_));
 OAI21_X1 _19764_ (.A(_03553_),
    .B1(_03558_),
    .B2(_03561_),
    .ZN(_03562_));
 NAND3_X2 _19765_ (.A1(_11070_),
    .A2(_11067_),
    .A3(_15860_),
    .ZN(_03563_));
 NOR2_X2 _19766_ (.A1(_15884_),
    .A2(_15892_),
    .ZN(_03564_));
 OAI21_X1 _19767_ (.A(_03564_),
    .B1(_03501_),
    .B2(_11066_),
    .ZN(_03565_));
 NOR2_X1 _19768_ (.A1(_15888_),
    .A2(_15892_),
    .ZN(_03566_));
 OAI221_X2 _19769_ (.A(_03566_),
    .B1(_03495_),
    .B2(_15860_),
    .C1(_03501_),
    .C2(_03503_),
    .ZN(_03567_));
 NOR3_X1 _19770_ (.A1(_10934_),
    .A2(_10975_),
    .A3(_03499_),
    .ZN(_03568_));
 OAI22_X2 _19771_ (.A1(_03563_),
    .A2(_03565_),
    .B1(_03567_),
    .B2(_03568_),
    .ZN(_03569_));
 NOR2_X1 _19772_ (.A1(_03495_),
    .A2(_15876_),
    .ZN(_03570_));
 AND3_X1 _19773_ (.A1(_15873_),
    .A2(_03570_),
    .A3(_03553_),
    .ZN(_03571_));
 AND3_X1 _19774_ (.A1(_11065_),
    .A2(_03570_),
    .A3(_03566_),
    .ZN(_03572_));
 AND2_X1 _19775_ (.A1(_03553_),
    .A2(_03572_),
    .ZN(_03573_));
 NOR3_X4 _19776_ (.A1(_03500_),
    .A2(_10744_),
    .A3(_03434_),
    .ZN(_03574_));
 NAND4_X4 _19777_ (.A1(_11070_),
    .A2(_11067_),
    .A3(_15860_),
    .A4(_03574_),
    .ZN(_03575_));
 OAI211_X4 _19778_ (.A(_03506_),
    .B(_15860_),
    .C1(_10975_),
    .C2(_10934_),
    .ZN(_03576_));
 NAND2_X2 _19779_ (.A1(_03506_),
    .A2(_03499_),
    .ZN(_03577_));
 NAND3_X1 _19780_ (.A1(_03575_),
    .A2(_03576_),
    .A3(_03577_),
    .ZN(_03578_));
 AOI22_X2 _19781_ (.A1(_03569_),
    .A2(_03571_),
    .B1(_03573_),
    .B2(_03578_),
    .ZN(_03579_));
 OAI211_X4 _19782_ (.A(_15860_),
    .B(_11065_),
    .C1(_10934_),
    .C2(_10975_),
    .ZN(_03580_));
 NAND2_X2 _19783_ (.A1(_15876_),
    .A2(_03574_),
    .ZN(_03581_));
 NOR3_X2 _19784_ (.A1(_03513_),
    .A2(_03580_),
    .A3(_03581_),
    .ZN(_03582_));
 AOI21_X1 _19785_ (.A(_03494_),
    .B1(_03564_),
    .B2(_03537_),
    .ZN(_03583_));
 AOI211_X2 _19786_ (.A(_03502_),
    .B(_03583_),
    .C1(_03539_),
    .C2(_10921_),
    .ZN(_03584_));
 OAI21_X1 _19787_ (.A(_03553_),
    .B1(_03582_),
    .B2(_03584_),
    .ZN(_03585_));
 NOR2_X1 _19788_ (.A1(_03495_),
    .A2(_03534_),
    .ZN(_03586_));
 NOR2_X2 _19789_ (.A1(_15892_),
    .A2(_15916_),
    .ZN(_03587_));
 AND4_X2 _19790_ (.A1(_15929_),
    .A2(_03491_),
    .A3(_03586_),
    .A4(_03587_),
    .ZN(_03588_));
 NOR3_X1 _19791_ (.A1(_03495_),
    .A2(_15880_),
    .A3(_03555_),
    .ZN(_03589_));
 OAI211_X2 _19792_ (.A(_03588_),
    .B(_03589_),
    .C1(_03506_),
    .C2(_03580_),
    .ZN(_03590_));
 AND2_X1 _19793_ (.A1(_03556_),
    .A2(_03535_),
    .ZN(_03591_));
 AND4_X1 _19794_ (.A1(_15869_),
    .A2(_03489_),
    .A3(_15929_),
    .A4(_03491_),
    .ZN(_03592_));
 OAI211_X2 _19795_ (.A(_11071_),
    .B(_03591_),
    .C1(_03592_),
    .C2(_03553_),
    .ZN(_03593_));
 NOR3_X4 _19796_ (.A1(_10934_),
    .A2(_10975_),
    .A3(_15864_),
    .ZN(_03594_));
 AND3_X2 _19797_ (.A1(_15869_),
    .A2(_03491_),
    .A3(_03485_),
    .ZN(_03595_));
 NAND3_X2 _19798_ (.A1(_11066_),
    .A2(_03493_),
    .A3(_11418_),
    .ZN(_03596_));
 NOR2_X1 _19799_ (.A1(_15876_),
    .A2(_03596_),
    .ZN(_03597_));
 NAND4_X1 _19800_ (.A1(_03564_),
    .A2(_03594_),
    .A3(_03595_),
    .A4(_03597_),
    .ZN(_03598_));
 AOI21_X1 _19801_ (.A(_15896_),
    .B1(_03502_),
    .B2(_03500_),
    .ZN(_03599_));
 AND3_X1 _19802_ (.A1(_15884_),
    .A2(_03570_),
    .A3(_03599_),
    .ZN(_03600_));
 NAND4_X1 _19803_ (.A1(_11065_),
    .A2(_11071_),
    .A3(_03492_),
    .A4(_03600_),
    .ZN(_03601_));
 AND4_X1 _19804_ (.A1(_03590_),
    .A2(_03593_),
    .A3(_03598_),
    .A4(_03601_),
    .ZN(_03602_));
 NAND4_X2 _19805_ (.A1(_03562_),
    .A2(_03579_),
    .A3(_03585_),
    .A4(_03602_),
    .ZN(_03603_));
 OAI21_X1 _19806_ (.A(_03509_),
    .B1(_03552_),
    .B2(_03603_),
    .ZN(_03604_));
 INV_X1 _19807_ (.A(_01161_),
    .ZN(_03605_));
 AOI21_X1 _19808_ (.A(_03480_),
    .B1(_03604_),
    .B2(_03605_),
    .ZN(_03606_));
 NOR2_X1 _19809_ (.A1(_03461_),
    .A2(_03606_),
    .ZN(\id_stage_i.controller_i.illegal_insn_d ));
 NOR2_X4 _19810_ (.A1(_10305_),
    .A2(_03435_),
    .ZN(_03607_));
 OR2_X2 _19811_ (.A1(_10891_),
    .A2(_10892_),
    .ZN(_03608_));
 NOR3_X4 _19812_ (.A1(_03467_),
    .A2(_03471_),
    .A3(_03608_),
    .ZN(_03609_));
 NOR2_X2 _19813_ (.A1(_03607_),
    .A2(_03609_),
    .ZN(_03610_));
 AOI21_X1 _19814_ (.A(_03461_),
    .B1(_03606_),
    .B2(_03610_),
    .ZN(\id_stage_i.controller_i.exc_req_d ));
 BUF_X4 _19815_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .Z(_03611_));
 NAND2_X4 _19816_ (.A1(_03611_),
    .A2(_03451_),
    .ZN(_03612_));
 CLKBUF_X3 _19817_ (.A(_03612_),
    .Z(_03613_));
 BUF_X4 _19818_ (.A(_03431_),
    .Z(_03614_));
 CLKBUF_X3 _19819_ (.A(_03441_),
    .Z(_03615_));
 OAI21_X1 _19820_ (.A(_03614_),
    .B1(_03615_),
    .B2(_03447_),
    .ZN(_03616_));
 NAND2_X1 _19821_ (.A1(_03613_),
    .A2(_03616_),
    .ZN(_00005_));
 BUF_X2 _19822_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Z(_03617_));
 NAND2_X1 _19823_ (.A1(_03617_),
    .A2(_03615_),
    .ZN(_03618_));
 BUF_X4 _19824_ (.A(_16105_),
    .Z(_03619_));
 INV_X2 _19825_ (.A(_03619_),
    .ZN(_03620_));
 XNOR2_X2 _19826_ (.A(_11735_),
    .B(_11726_),
    .ZN(\alu_adder_result_ex[5] ));
 OAI21_X1 _19827_ (.A(_11841_),
    .B1(_11719_),
    .B2(_11842_),
    .ZN(_03621_));
 XOR2_X2 _19828_ (.A(_11721_),
    .B(_03621_),
    .Z(\alu_adder_result_ex[3] ));
 OR3_X1 _19829_ (.A1(_03620_),
    .A2(\alu_adder_result_ex[5] ),
    .A3(\alu_adder_result_ex[3] ),
    .ZN(_03622_));
 OR4_X1 _19830_ (.A1(\alu_adder_result_ex[7] ),
    .A2(\alu_adder_result_ex[9] ),
    .A3(\alu_adder_result_ex[11] ),
    .A4(_03622_),
    .ZN(_03623_));
 OR3_X1 _19831_ (.A1(\alu_adder_result_ex[13] ),
    .A2(\alu_adder_result_ex[15] ),
    .A3(_03623_),
    .ZN(_03624_));
 OR3_X1 _19832_ (.A1(\alu_adder_result_ex[6] ),
    .A2(\alu_adder_result_ex[8] ),
    .A3(_03624_),
    .ZN(_03625_));
 OR2_X1 _19833_ (.A1(\alu_adder_result_ex[17] ),
    .A2(\alu_adder_result_ex[21] ),
    .ZN(_03626_));
 OR4_X2 _19834_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_12101_),
    .A3(_03625_),
    .A4(_03626_),
    .ZN(_03627_));
 INV_X1 _19835_ (.A(_11744_),
    .ZN(_03628_));
 AOI221_X2 _19836_ (.A(_15371_),
    .B1(_14064_),
    .B2(_03628_),
    .C1(_15373_),
    .C2(_10815_),
    .ZN(_03629_));
 XNOR2_X2 _19837_ (.A(_11720_),
    .B(_03629_),
    .ZN(\alu_adder_result_ex[2] ));
 NOR2_X1 _19838_ (.A1(_11722_),
    .A2(_11838_),
    .ZN(_03630_));
 MUX2_X1 _19839_ (.A(_11722_),
    .B(_03630_),
    .S(_11844_),
    .Z(_03631_));
 NAND2_X1 _19840_ (.A1(_11722_),
    .A2(_11838_),
    .ZN(_03632_));
 NOR2_X1 _19841_ (.A1(_11401_),
    .A2(_11862_),
    .ZN(_03633_));
 AOI211_X2 _19842_ (.A(_11854_),
    .B(_03632_),
    .C1(_03633_),
    .C2(_11858_),
    .ZN(_03634_));
 AND2_X1 _19843_ (.A1(_11725_),
    .A2(_11844_),
    .ZN(_03635_));
 AOI211_X4 _19844_ (.A(_03631_),
    .B(_03634_),
    .C1(_03635_),
    .C2(_11514_),
    .ZN(\alu_adder_result_ex[4] ));
 OR2_X1 _19845_ (.A1(\alu_adder_result_ex[19] ),
    .A2(\alu_adder_result_ex[4] ),
    .ZN(_03636_));
 OR4_X2 _19846_ (.A1(\alu_adder_result_ex[16] ),
    .A2(\alu_adder_result_ex[23] ),
    .A3(\alu_adder_result_ex[2] ),
    .A4(_03636_),
    .ZN(_03637_));
 NAND2_X1 _19847_ (.A1(_12593_),
    .A2(_13111_),
    .ZN(_03638_));
 NAND2_X1 _19848_ (.A1(_12594_),
    .A2(_13111_),
    .ZN(_03639_));
 MUX2_X1 _19849_ (.A(_03638_),
    .B(_03639_),
    .S(_12610_),
    .Z(_03640_));
 OR2_X1 _19850_ (.A1(\alu_adder_result_ex[27] ),
    .A2(net14),
    .ZN(_03641_));
 OR4_X2 _19851_ (.A1(\alu_adder_result_ex[14] ),
    .A2(net382),
    .A3(_03640_),
    .A4(_03641_),
    .ZN(_03642_));
 OR4_X4 _19852_ (.A1(_03430_),
    .A2(_03627_),
    .A3(_03637_),
    .A4(_03642_),
    .ZN(_03643_));
 OR2_X1 _19853_ (.A1(\alu_adder_result_ex[20] ),
    .A2(\alu_adder_result_ex[28] ),
    .ZN(_03644_));
 OR4_X2 _19854_ (.A1(\alu_adder_result_ex[22] ),
    .A2(\alu_adder_result_ex[24] ),
    .A3(\alu_adder_result_ex[31] ),
    .A4(_03644_),
    .ZN(_03645_));
 NOR2_X2 _19855_ (.A1(_03643_),
    .A2(_03645_),
    .ZN(_03646_));
 CLKBUF_X3 _19856_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .Z(_03647_));
 NAND2_X1 _19857_ (.A1(_03647_),
    .A2(_03451_),
    .ZN(_03648_));
 OAI21_X1 _19858_ (.A(_03618_),
    .B1(_03646_),
    .B2(_03648_),
    .ZN(_00004_));
 NAND2_X1 _19859_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .A2(_03615_),
    .ZN(_03649_));
 BUF_X4 _19860_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Z(_03650_));
 BUF_X4 _19861_ (.A(_03650_),
    .Z(_03651_));
 BUF_X4 _19862_ (.A(_03651_),
    .Z(_03652_));
 AOI21_X1 _19863_ (.A(_03652_),
    .B1(_03647_),
    .B2(_03646_),
    .ZN(_03653_));
 OAI21_X1 _19864_ (.A(_03649_),
    .B1(_03653_),
    .B2(_03615_),
    .ZN(_00003_));
 INV_X4 _19865_ (.A(_14068_),
    .ZN(\alu_adder_result_ex[0] ));
 OR2_X1 _19866_ (.A1(_11430_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .ZN(_03654_));
 CLKBUF_X3 _19867_ (.A(_03654_),
    .Z(_03655_));
 BUF_X4 _19868_ (.A(_03655_),
    .Z(_03656_));
 NAND2_X4 _19869_ (.A1(_12316_),
    .A2(_03656_),
    .ZN(_03657_));
 BUF_X4 _19870_ (.A(_03656_),
    .Z(_03658_));
 OR2_X1 _19871_ (.A1(_10706_),
    .A2(_10729_),
    .ZN(_03659_));
 BUF_X4 _19872_ (.A(_03659_),
    .Z(_03660_));
 OAI21_X4 _19873_ (.A(_03657_),
    .B1(_03658_),
    .B2(_03660_),
    .ZN(_03661_));
 INV_X4 _19874_ (.A(_03661_),
    .ZN(_03662_));
 OR2_X2 _19875_ (.A1(_11400_),
    .A2(_11430_),
    .ZN(_03663_));
 BUF_X4 _19876_ (.A(_03663_),
    .Z(_03664_));
 NOR2_X1 _19877_ (.A1(net411),
    .A2(_03664_),
    .ZN(_03665_));
 BUF_X4 _19878_ (.A(_03663_),
    .Z(_03666_));
 AOI21_X4 _19879_ (.A(_03665_),
    .B1(_03666_),
    .B2(_12350_),
    .ZN(_03667_));
 NOR2_X1 _19880_ (.A1(_03662_),
    .A2(_03667_),
    .ZN(_15550_));
 OR2_X1 _19881_ (.A1(_00217_),
    .A2(_11402_),
    .ZN(_03668_));
 CLKBUF_X3 _19882_ (.A(_11433_),
    .Z(_03669_));
 BUF_X2 _19883_ (.A(_00690_),
    .Z(_03670_));
 OAI21_X1 _19884_ (.A(_03668_),
    .B1(_03669_),
    .B2(_03670_),
    .ZN(_03671_));
 AOI22_X1 _19885_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A2(_03658_),
    .B1(_03671_),
    .B2(_11431_),
    .ZN(_03672_));
 INV_X1 _19886_ (.A(_03672_),
    .ZN(_15551_));
 INV_X2 _19887_ (.A(_03667_),
    .ZN(_03673_));
 AND2_X2 _19888_ (.A1(_11928_),
    .A2(_10433_),
    .ZN(_03674_));
 AOI21_X4 _19889_ (.A(_03674_),
    .B1(_10470_),
    .B2(_10474_),
    .ZN(_03675_));
 MUX2_X2 _19890_ (.A(_03675_),
    .B(_12392_),
    .S(_03656_),
    .Z(_03676_));
 NAND2_X1 _19891_ (.A1(_03673_),
    .A2(net339),
    .ZN(_14069_));
 BUF_X4 _19892_ (.A(_03667_),
    .Z(_03677_));
 NOR2_X1 _19893_ (.A1(_10972_),
    .A2(_03655_),
    .ZN(_03678_));
 AOI21_X4 _19894_ (.A(_03678_),
    .B1(_03656_),
    .B2(net346),
    .ZN(_03679_));
 NOR2_X1 _19895_ (.A1(_03677_),
    .A2(_03679_),
    .ZN(_15563_));
 BUF_X8 _19896_ (.A(_03676_),
    .Z(_03680_));
 AND2_X2 _19897_ (.A1(_10642_),
    .A2(_10659_),
    .ZN(_03681_));
 MUX2_X1 _19898_ (.A(_03681_),
    .B(_12425_),
    .S(_03663_),
    .Z(_03682_));
 BUF_X4 _19899_ (.A(_03682_),
    .Z(_03683_));
 NAND2_X1 _19900_ (.A1(net338),
    .A2(_03683_),
    .ZN(_14076_));
 AND2_X4 _19901_ (.A1(net349),
    .A2(_03655_),
    .ZN(_03684_));
 NOR2_X4 _19902_ (.A1(_11430_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .ZN(_03685_));
 AOI21_X4 _19903_ (.A(_03684_),
    .B1(_03685_),
    .B2(_11019_),
    .ZN(_03686_));
 NOR2_X1 _19904_ (.A1(_03677_),
    .A2(_03686_),
    .ZN(_15567_));
 BUF_X4 _19905_ (.A(_03679_),
    .Z(_03687_));
 INV_X2 _19906_ (.A(_03683_),
    .ZN(_03688_));
 NOR2_X1 _19907_ (.A1(_03687_),
    .A2(_03688_),
    .ZN(_15566_));
 MUX2_X1 _19908_ (.A(net293),
    .B(_12514_),
    .S(_03666_),
    .Z(_03689_));
 BUF_X4 _19909_ (.A(_03689_),
    .Z(_03690_));
 NAND2_X1 _19910_ (.A1(net338),
    .A2(_03690_),
    .ZN(_14080_));
 NOR2_X1 _19911_ (.A1(_11057_),
    .A2(_03656_),
    .ZN(_03691_));
 AOI21_X4 _19912_ (.A(_03691_),
    .B1(_03656_),
    .B2(_12651_),
    .ZN(_03692_));
 NOR2_X1 _19913_ (.A1(_03677_),
    .A2(_03692_),
    .ZN(_14084_));
 NOR2_X1 _19914_ (.A1(_03688_),
    .A2(_03686_),
    .ZN(_14086_));
 INV_X2 _19915_ (.A(_03689_),
    .ZN(_03693_));
 NOR2_X1 _19916_ (.A1(_03687_),
    .A2(_03693_),
    .ZN(_14085_));
 MUX2_X2 _19917_ (.A(net319),
    .B(_12589_),
    .S(_03664_),
    .Z(_03694_));
 BUF_X4 _19918_ (.A(_03694_),
    .Z(_03695_));
 NAND2_X1 _19919_ (.A1(net338),
    .A2(_03695_),
    .ZN(_14091_));
 NAND4_X4 _19920_ (.A1(_11083_),
    .A2(_11093_),
    .A3(_11105_),
    .A4(_11114_),
    .ZN(_03696_));
 MUX2_X2 _19921_ (.A(_03696_),
    .B(_12725_),
    .S(_03656_),
    .Z(_03697_));
 INV_X1 _19922_ (.A(_03697_),
    .ZN(_03698_));
 NOR2_X1 _19923_ (.A1(_03677_),
    .A2(_03698_),
    .ZN(_15589_));
 NOR2_X1 _19924_ (.A1(_03688_),
    .A2(_03692_),
    .ZN(_14105_));
 BUF_X8 _19925_ (.A(_03686_),
    .Z(_03699_));
 NOR2_X1 _19926_ (.A1(_03699_),
    .A2(_03693_),
    .ZN(_14104_));
 INV_X2 _19927_ (.A(_03694_),
    .ZN(_03700_));
 NOR2_X1 _19928_ (.A1(_03687_),
    .A2(_03700_),
    .ZN(_14106_));
 MUX2_X2 _19929_ (.A(_11591_),
    .B(net358),
    .S(_03666_),
    .Z(_03701_));
 BUF_X4 _19930_ (.A(_03701_),
    .Z(_03702_));
 NAND2_X1 _19931_ (.A1(net338),
    .A2(_03702_),
    .ZN(_14110_));
 MUX2_X2 _19932_ (.A(_11158_),
    .B(_12823_),
    .S(_03655_),
    .Z(_03703_));
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 INV_X1 _19934_ (.A(net324),
    .ZN(_03705_));
 NOR2_X1 _19935_ (.A1(_03677_),
    .A2(_03705_),
    .ZN(_15602_));
 NOR2_X1 _19936_ (.A1(_03688_),
    .A2(_03698_),
    .ZN(_15601_));
 NOR2_X1 _19937_ (.A1(_03693_),
    .A2(_03692_),
    .ZN(_14127_));
 NOR2_X1 _19938_ (.A1(_03699_),
    .A2(_03700_),
    .ZN(_14129_));
 INV_X2 _19939_ (.A(_03701_),
    .ZN(_03706_));
 NOR2_X1 _19940_ (.A1(_03687_),
    .A2(_03706_),
    .ZN(_14128_));
 MUX2_X1 _19941_ (.A(_11629_),
    .B(net361),
    .S(_03666_),
    .Z(_03707_));
 BUF_X4 _19942_ (.A(_03707_),
    .Z(_03708_));
 NAND2_X1 _19943_ (.A1(net338),
    .A2(_03708_),
    .ZN(_14132_));
 MUX2_X2 _19944_ (.A(_11202_),
    .B(net421),
    .S(_03655_),
    .Z(_03709_));
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 NAND2_X1 _19946_ (.A1(_03673_),
    .A2(net322),
    .ZN(_14146_));
 CLKBUF_X3 _19947_ (.A(_03692_),
    .Z(_03711_));
 NOR2_X1 _19948_ (.A1(_03711_),
    .A2(_03700_),
    .ZN(_14152_));
 NOR2_X1 _19949_ (.A1(_03699_),
    .A2(_03706_),
    .ZN(_14151_));
 INV_X2 _19950_ (.A(_03707_),
    .ZN(_03712_));
 NOR2_X1 _19951_ (.A1(_03687_),
    .A2(_03712_),
    .ZN(_14150_));
 NOR2_X4 _19952_ (.A1(_12840_),
    .A2(_12858_),
    .ZN(_03713_));
 MUX2_X1 _19953_ (.A(_11672_),
    .B(_03713_),
    .S(_03666_),
    .Z(_03714_));
 BUF_X4 _19954_ (.A(_03714_),
    .Z(_03715_));
 NAND2_X1 _19955_ (.A1(_03680_),
    .A2(_03715_),
    .ZN(_14161_));
 NAND2_X4 _19956_ (.A1(_12985_),
    .A2(_03656_),
    .ZN(_03716_));
 OAI21_X4 _19957_ (.A(_03716_),
    .B1(_03658_),
    .B2(_11241_),
    .ZN(_03717_));
 INV_X1 _19958_ (.A(net336),
    .ZN(_03718_));
 NOR2_X1 _19959_ (.A1(_03677_),
    .A2(_03718_),
    .ZN(_15635_));
 NAND2_X1 _19960_ (.A1(_03683_),
    .A2(net322),
    .ZN(_14178_));
 NOR2_X1 _19961_ (.A1(_03711_),
    .A2(_03706_),
    .ZN(_14183_));
 NOR2_X1 _19962_ (.A1(_03699_),
    .A2(_03712_),
    .ZN(_14182_));
 NOR2_X2 _19963_ (.A1(_11431_),
    .A2(_11430_),
    .ZN(_03719_));
 BUF_X4 _19964_ (.A(_03719_),
    .Z(_03720_));
 NOR2_X1 _19965_ (.A1(_12859_),
    .A2(_03720_),
    .ZN(_03721_));
 AOI21_X4 _19966_ (.A(_03721_),
    .B1(_03720_),
    .B2(_11672_),
    .ZN(_03722_));
 NOR2_X1 _19967_ (.A1(_03687_),
    .A2(_03722_),
    .ZN(_14184_));
 NOR2_X4 _19968_ (.A1(_11694_),
    .A2(_11713_),
    .ZN(_03723_));
 NOR2_X4 _19969_ (.A1(_12915_),
    .A2(_12933_),
    .ZN(_03724_));
 MUX2_X1 _19970_ (.A(_03723_),
    .B(_03724_),
    .S(_03666_),
    .Z(_03725_));
 BUF_X4 _19971_ (.A(_03725_),
    .Z(_03726_));
 NAND2_X1 _19972_ (.A1(_03680_),
    .A2(_03726_),
    .ZN(_14190_));
 OR4_X4 _19973_ (.A1(_11253_),
    .A2(_11260_),
    .A3(_11269_),
    .A4(_11278_),
    .ZN(_03727_));
 MUX2_X1 _19974_ (.A(_03727_),
    .B(_13061_),
    .S(_03655_),
    .Z(_03728_));
 BUF_X4 _19975_ (.A(_03728_),
    .Z(_03729_));
 INV_X1 _19976_ (.A(_03729_),
    .ZN(_03730_));
 NOR2_X1 _19977_ (.A1(_03677_),
    .A2(_03730_),
    .ZN(_15645_));
 NOR2_X1 _19978_ (.A1(_03688_),
    .A2(_03718_),
    .ZN(_15646_));
 NAND2_X1 _19979_ (.A1(_03690_),
    .A2(_03709_),
    .ZN(_14208_));
 NOR2_X1 _19980_ (.A1(_03711_),
    .A2(_03712_),
    .ZN(_14215_));
 NOR2_X2 _19981_ (.A1(_03699_),
    .A2(_03722_),
    .ZN(_14214_));
 MUX2_X2 _19982_ (.A(_11714_),
    .B(_12934_),
    .S(_03666_),
    .Z(_03731_));
 NOR2_X1 _19983_ (.A1(_03687_),
    .A2(_03731_),
    .ZN(_14213_));
 NOR2_X4 _19984_ (.A1(_11764_),
    .A2(_11786_),
    .ZN(_03732_));
 NOR2_X4 _19985_ (.A1(_13004_),
    .A2(_13022_),
    .ZN(_03733_));
 MUX2_X1 _19986_ (.A(_03732_),
    .B(_03733_),
    .S(_03666_),
    .Z(_03734_));
 BUF_X4 _19987_ (.A(_03734_),
    .Z(_03735_));
 NAND2_X1 _19988_ (.A1(_03680_),
    .A2(_03735_),
    .ZN(_14221_));
 AND2_X2 _19989_ (.A1(_11296_),
    .A2(_11312_),
    .ZN(_03736_));
 MUX2_X1 _19990_ (.A(_03736_),
    .B(_13155_),
    .S(_03655_),
    .Z(_03737_));
 BUF_X4 _19991_ (.A(_03737_),
    .Z(_03738_));
 BUF_X4 _19992_ (.A(_03738_),
    .Z(_03739_));
 NAND2_X1 _19993_ (.A1(_03673_),
    .A2(_03739_),
    .ZN(_14243_));
 NAND2_X1 _19994_ (.A1(_03695_),
    .A2(_03709_),
    .ZN(_14248_));
 NOR2_X1 _19995_ (.A1(_03711_),
    .A2(_03722_),
    .ZN(_14255_));
 NOR2_X2 _19996_ (.A1(_03699_),
    .A2(_03731_),
    .ZN(_14254_));
 MUX2_X2 _19997_ (.A(_11787_),
    .B(_13023_),
    .S(_03666_),
    .Z(_03740_));
 NOR2_X2 _19998_ (.A1(_03687_),
    .A2(_03740_),
    .ZN(_14253_));
 MUX2_X1 _19999_ (.A(_11824_),
    .B(_13097_),
    .S(_03666_),
    .Z(_03741_));
 BUF_X4 _20000_ (.A(_03741_),
    .Z(_03742_));
 NAND2_X1 _20001_ (.A1(_03680_),
    .A2(_03742_),
    .ZN(_14261_));
 NOR4_X4 _20002_ (.A1(_11328_),
    .A2(_11335_),
    .A3(_11342_),
    .A4(_11350_),
    .ZN(_03743_));
 NOR2_X1 _20003_ (.A1(_03743_),
    .A2(_03655_),
    .ZN(_03744_));
 AOI21_X4 _20004_ (.A(_03744_),
    .B1(_03656_),
    .B2(_13224_),
    .ZN(_03745_));
 CLKBUF_X3 _20005_ (.A(_03745_),
    .Z(_03746_));
 NOR2_X1 _20006_ (.A1(_03677_),
    .A2(_03746_),
    .ZN(_15677_));
 NAND2_X1 _20007_ (.A1(_03683_),
    .A2(_03739_),
    .ZN(_14283_));
 NAND2_X1 _20008_ (.A1(_03702_),
    .A2(_03709_),
    .ZN(_14288_));
 NOR2_X1 _20009_ (.A1(_03711_),
    .A2(_03731_),
    .ZN(_14295_));
 NOR2_X2 _20010_ (.A1(_03699_),
    .A2(_03740_),
    .ZN(_14294_));
 NOR3_X2 _20011_ (.A1(_13078_),
    .A2(_13096_),
    .A3(_03720_),
    .ZN(_03747_));
 AOI21_X4 _20012_ (.A(_03747_),
    .B1(_03720_),
    .B2(_11824_),
    .ZN(_03748_));
 NOR2_X2 _20013_ (.A1(_03687_),
    .A2(_03748_),
    .ZN(_14293_));
 MUX2_X2 _20014_ (.A(_11898_),
    .B(net350),
    .S(_03664_),
    .Z(_03749_));
 NOR2_X2 clone93 (.A1(_03780_),
    .A2(_03685_),
    .ZN(net364));
 NAND2_X4 _20016_ (.A1(_03680_),
    .A2(_03749_),
    .ZN(_14304_));
 AND2_X1 _20017_ (.A1(_11993_),
    .A2(_03685_),
    .ZN(_03751_));
 AOI21_X2 _20018_ (.A(_03751_),
    .B1(_03656_),
    .B2(_13314_),
    .ZN(_03752_));
 CLKBUF_X3 _20019_ (.A(_03752_),
    .Z(_03753_));
 NOR2_X1 _20020_ (.A1(_03677_),
    .A2(_03753_),
    .ZN(_15688_));
 NOR2_X1 _20021_ (.A1(_03688_),
    .A2(_03746_),
    .ZN(_15687_));
 NAND2_X1 _20022_ (.A1(_03690_),
    .A2(_03739_),
    .ZN(_14327_));
 NAND2_X1 _20023_ (.A1(_03708_),
    .A2(_03709_),
    .ZN(_14331_));
 NOR2_X1 _20024_ (.A1(_03711_),
    .A2(_03740_),
    .ZN(_14338_));
 NOR2_X2 _20025_ (.A1(_03699_),
    .A2(_03748_),
    .ZN(_14337_));
 INV_X2 _20026_ (.A(_03749_),
    .ZN(_03754_));
 NOR2_X2 _20027_ (.A1(_03687_),
    .A2(_03754_),
    .ZN(_14336_));
 MUX2_X2 _20028_ (.A(net365),
    .B(net340),
    .S(_03664_),
    .Z(_03755_));
 BUF_X4 _20029_ (.A(_03755_),
    .Z(_03756_));
 NAND2_X1 _20030_ (.A1(net339),
    .A2(_03756_),
    .ZN(_14354_));
 AND2_X2 _20031_ (.A1(_12044_),
    .A2(_03685_),
    .ZN(_03757_));
 AOI21_X2 _20032_ (.A(_03757_),
    .B1(_03658_),
    .B2(_03166_),
    .ZN(_03758_));
 BUF_X4 _20033_ (.A(_03758_),
    .Z(_03759_));
 NOR2_X1 _20034_ (.A1(_03667_),
    .A2(_03759_),
    .ZN(_14374_));
 NOR2_X1 _20035_ (.A1(_03688_),
    .A2(_03753_),
    .ZN(_14373_));
 NOR2_X1 _20036_ (.A1(_03693_),
    .A2(_03746_),
    .ZN(_14372_));
 NAND2_X1 _20037_ (.A1(_03695_),
    .A2(_03738_),
    .ZN(_14377_));
 BUF_X8 _20038_ (.A(_03709_),
    .Z(_03760_));
 NAND2_X1 _20039_ (.A1(_03760_),
    .A2(_03715_),
    .ZN(_14386_));
 NOR2_X1 _20040_ (.A1(_03711_),
    .A2(_03748_),
    .ZN(_14390_));
 NOR2_X1 _20041_ (.A1(_03699_),
    .A2(_03754_),
    .ZN(_14392_));
 INV_X2 _20042_ (.A(_03755_),
    .ZN(_03761_));
 NOR2_X1 _20043_ (.A1(_03679_),
    .A2(_03761_),
    .ZN(_14391_));
 OR2_X4 _20044_ (.A1(_03112_),
    .A2(_03130_),
    .ZN(_03762_));
 MUX2_X2 _20045_ (.A(_10868_),
    .B(_03762_),
    .S(_03664_),
    .Z(_03763_));
 CLKBUF_X3 _20046_ (.A(_03763_),
    .Z(_03764_));
 NAND2_X1 _20047_ (.A1(net339),
    .A2(_03764_),
    .ZN(_14406_));
 MUX2_X2 _20048_ (.A(_12144_),
    .B(_03275_),
    .S(_03655_),
    .Z(_03765_));
 INV_X1 _20049_ (.A(_03765_),
    .ZN(_03766_));
 NOR2_X1 _20050_ (.A1(_03667_),
    .A2(_03766_),
    .ZN(_15708_));
 INV_X2 _20051_ (.A(_03758_),
    .ZN(_03767_));
 NAND2_X1 _20052_ (.A1(_03683_),
    .A2(_03767_),
    .ZN(_14430_));
 NAND2_X1 _20053_ (.A1(_03702_),
    .A2(_03738_),
    .ZN(_14434_));
 NAND2_X4 _20054_ (.A1(_03760_),
    .A2(_03726_),
    .ZN(_14442_));
 NOR2_X1 _20055_ (.A1(_03711_),
    .A2(_03754_),
    .ZN(_14446_));
 NOR2_X2 _20056_ (.A1(_03699_),
    .A2(_03761_),
    .ZN(_14448_));
 INV_X1 _20057_ (.A(_03763_),
    .ZN(_03768_));
 NOR2_X1 _20058_ (.A1(_03679_),
    .A2(_03768_),
    .ZN(_14447_));
 OR2_X4 _20059_ (.A1(_03185_),
    .A2(_03203_),
    .ZN(_03769_));
 MUX2_X2 _20060_ (.A(_12075_),
    .B(_03769_),
    .S(_03664_),
    .Z(_03770_));
 CLKBUF_X3 _20061_ (.A(_03770_),
    .Z(_03771_));
 NAND2_X1 _20062_ (.A1(net339),
    .A2(_03771_),
    .ZN(_14461_));
 INV_X2 _20063_ (.A(_03400_),
    .ZN(_03772_));
 MUX2_X1 _20064_ (.A(net327),
    .B(_03772_),
    .S(_03655_),
    .Z(_03773_));
 BUF_X4 _20065_ (.A(_03773_),
    .Z(_03774_));
 AND2_X1 _20066_ (.A1(_03673_),
    .A2(_03774_),
    .ZN(_15719_));
 NOR2_X1 _20067_ (.A1(_03688_),
    .A2(_03766_),
    .ZN(_15718_));
 NOR2_X1 _20068_ (.A1(_03693_),
    .A2(_03759_),
    .ZN(_14484_));
 NOR2_X1 _20069_ (.A1(_03700_),
    .A2(_03753_),
    .ZN(_14483_));
 NOR2_X1 _20070_ (.A1(_03706_),
    .A2(_03746_),
    .ZN(_14482_));
 NAND2_X1 _20071_ (.A1(_03708_),
    .A2(_03738_),
    .ZN(_14489_));
 NAND2_X2 _20072_ (.A1(_03760_),
    .A2(_03735_),
    .ZN(_14500_));
 NOR2_X1 _20073_ (.A1(_03711_),
    .A2(_03761_),
    .ZN(_14505_));
 NOR2_X1 _20074_ (.A1(_03686_),
    .A2(_03768_),
    .ZN(_14504_));
 INV_X1 _20075_ (.A(_03770_),
    .ZN(_03775_));
 NOR2_X1 _20076_ (.A1(_03679_),
    .A2(_03775_),
    .ZN(_14506_));
 MUX2_X2 _20077_ (.A(_12177_),
    .B(_03311_),
    .S(_03664_),
    .Z(_03776_));
 CLKBUF_X3 _20078_ (.A(_03776_),
    .Z(_03777_));
 NAND2_X1 _20079_ (.A1(_03676_),
    .A2(_03777_),
    .ZN(_14520_));
 OR3_X1 _20080_ (.A1(_10550_),
    .A2(_11405_),
    .A3(_03400_),
    .ZN(_03778_));
 CLKBUF_X3 _20081_ (.A(_03778_),
    .Z(_03779_));
 BUF_X4 _20082_ (.A(_03779_),
    .Z(_03780_));
 NOR2_X4 _20083_ (.A1(_03780_),
    .A2(_03685_),
    .ZN(_03781_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 NAND2_X1 _20085_ (.A1(_03677_),
    .A2(_03781_),
    .ZN(_14539_));
 NOR2_X1 _20086_ (.A1(_03700_),
    .A2(_03759_),
    .ZN(_14545_));
 NOR2_X1 _20087_ (.A1(_03706_),
    .A2(_03753_),
    .ZN(_14544_));
 NOR2_X1 _20088_ (.A1(_03712_),
    .A2(_03746_),
    .ZN(_14546_));
 NAND2_X1 _20089_ (.A1(_03715_),
    .A2(_03738_),
    .ZN(_14554_));
 NAND2_X1 _20090_ (.A1(_03760_),
    .A2(_03742_),
    .ZN(_14565_));
 NOR2_X1 _20091_ (.A1(_03711_),
    .A2(_03768_),
    .ZN(_14572_));
 NOR2_X1 _20092_ (.A1(_03686_),
    .A2(_03775_),
    .ZN(_14571_));
 INV_X1 _20093_ (.A(_03776_),
    .ZN(_03782_));
 NOR2_X1 _20094_ (.A1(_03679_),
    .A2(_03782_),
    .ZN(_14570_));
 OR2_X2 _20095_ (.A1(_03371_),
    .A2(_03386_),
    .ZN(_03783_));
 MUX2_X2 _20096_ (.A(_12254_),
    .B(_03783_),
    .S(_03664_),
    .Z(_03784_));
 AND2_X1 _20097_ (.A1(_03676_),
    .A2(_03784_),
    .ZN(_14584_));
 BUF_X2 _20098_ (.A(_03664_),
    .Z(_03785_));
 INV_X1 _20099_ (.A(_03783_),
    .ZN(_03786_));
 NOR4_X2 _20100_ (.A1(_10310_),
    .A2(_10488_),
    .A3(_10346_),
    .A4(_10874_),
    .ZN(_03787_));
 AOI21_X2 _20101_ (.A(_10381_),
    .B1(_10380_),
    .B2(_10402_),
    .ZN(_03788_));
 OAI21_X4 _20102_ (.A(_11401_),
    .B1(_03787_),
    .B2(_03788_),
    .ZN(_03789_));
 NOR2_X4 _20103_ (.A1(_03786_),
    .A2(_03789_),
    .ZN(_03790_));
 BUF_X4 _20104_ (.A(_03790_),
    .Z(_03791_));
 NAND2_X4 _20105_ (.A1(_03785_),
    .A2(_03791_),
    .ZN(_03792_));
 NOR2_X4 _20106_ (.A1(_03792_),
    .A2(_03662_),
    .ZN(_14586_));
 NAND2_X1 _20107_ (.A1(_11430_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .ZN(_03793_));
 NAND2_X1 _20108_ (.A1(_11400_),
    .A2(_11433_),
    .ZN(_03794_));
 CLKBUF_X3 _20109_ (.A(_03794_),
    .Z(_03795_));
 OAI21_X1 _20110_ (.A(_03793_),
    .B1(_03795_),
    .B2(_03670_),
    .ZN(_14585_));
 NAND2_X1 _20111_ (.A1(_03688_),
    .A2(_03781_),
    .ZN(_14610_));
 NOR2_X1 _20112_ (.A1(_03706_),
    .A2(_03759_),
    .ZN(_14614_));
 NOR2_X1 _20113_ (.A1(_03712_),
    .A2(_03753_),
    .ZN(_14616_));
 NOR2_X1 _20114_ (.A1(_03722_),
    .A2(_03746_),
    .ZN(_14615_));
 NAND2_X1 _20115_ (.A1(_03726_),
    .A2(_03738_),
    .ZN(_14624_));
 NAND2_X1 _20116_ (.A1(_03760_),
    .A2(_03749_),
    .ZN(_14634_));
 NOR2_X1 _20117_ (.A1(_03692_),
    .A2(_03775_),
    .ZN(_14638_));
 NOR2_X1 _20118_ (.A1(_03686_),
    .A2(_03782_),
    .ZN(_14640_));
 INV_X1 _20119_ (.A(_03784_),
    .ZN(_03796_));
 NOR2_X1 _20120_ (.A1(_03679_),
    .A2(_03796_),
    .ZN(_14639_));
 NOR3_X2 _20121_ (.A1(_03786_),
    .A2(_03719_),
    .A3(_03789_),
    .ZN(_03797_));
 BUF_X4 _20122_ (.A(_03797_),
    .Z(_03798_));
 AND2_X4 _20123_ (.A1(_03676_),
    .A2(_03798_),
    .ZN(_14651_));
 NAND2_X1 _20124_ (.A1(_11430_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .ZN(_03799_));
 BUF_X2 _20125_ (.A(_00721_),
    .Z(_03800_));
 OAI21_X1 _20126_ (.A(_03799_),
    .B1(_03795_),
    .B2(_03800_),
    .ZN(_14652_));
 NAND2_X1 _20127_ (.A1(_03693_),
    .A2(_03781_),
    .ZN(_14671_));
 NOR2_X1 _20128_ (.A1(_03712_),
    .A2(_03759_),
    .ZN(_14675_));
 NOR2_X1 _20129_ (.A1(_03722_),
    .A2(_03753_),
    .ZN(_14674_));
 NOR2_X1 _20130_ (.A1(_03731_),
    .A2(_03746_),
    .ZN(_14676_));
 NAND2_X1 _20131_ (.A1(_03735_),
    .A2(_03738_),
    .ZN(_14683_));
 NAND2_X1 _20132_ (.A1(net321),
    .A2(_03756_),
    .ZN(_14694_));
 NOR2_X1 _20133_ (.A1(_03692_),
    .A2(_03782_),
    .ZN(_14698_));
 NOR2_X1 _20134_ (.A1(_03686_),
    .A2(_03796_),
    .ZN(_14697_));
 OR2_X1 _20135_ (.A1(_03679_),
    .A2(_03792_),
    .ZN(_14757_));
 INV_X1 _20136_ (.A(_14757_),
    .ZN(_14699_));
 OR3_X1 _20137_ (.A1(_00555_),
    .A2(_00132_),
    .A3(_03789_),
    .ZN(_03801_));
 BUF_X2 _20138_ (.A(_03801_),
    .Z(_03802_));
 CLKBUF_X3 _20139_ (.A(_03802_),
    .Z(_03803_));
 BUF_X2 _20140_ (.A(_00752_),
    .Z(_03804_));
 OAI21_X1 _20141_ (.A(_03803_),
    .B1(_03795_),
    .B2(_03804_),
    .ZN(_03805_));
 AND2_X1 _20142_ (.A1(_03785_),
    .A2(_03805_),
    .ZN(_14709_));
 NAND2_X1 _20143_ (.A1(_03700_),
    .A2(_03781_),
    .ZN(_14729_));
 NOR2_X1 _20144_ (.A1(_03722_),
    .A2(_03759_),
    .ZN(_14733_));
 NOR2_X1 _20145_ (.A1(_03731_),
    .A2(_03753_),
    .ZN(_14732_));
 NOR2_X1 _20146_ (.A1(_03740_),
    .A2(_03746_),
    .ZN(_14734_));
 NAND2_X1 _20147_ (.A1(_03739_),
    .A2(_03742_),
    .ZN(_14741_));
 NAND2_X1 _20148_ (.A1(net321),
    .A2(_03764_),
    .ZN(_14752_));
 OR2_X1 _20149_ (.A1(_03692_),
    .A2(_03796_),
    .ZN(_14756_));
 OR2_X1 _20150_ (.A1(_03686_),
    .A2(_03792_),
    .ZN(_14755_));
 INV_X1 _20151_ (.A(_14755_),
    .ZN(_14814_));
 INV_X2 _20152_ (.A(_00783_),
    .ZN(_03806_));
 NAND2_X1 _20153_ (.A1(_03806_),
    .A2(_11434_),
    .ZN(_03807_));
 AOI21_X1 _20154_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03807_),
    .ZN(_14766_));
 NAND2_X1 _20155_ (.A1(_03706_),
    .A2(_03781_),
    .ZN(_14786_));
 NOR2_X1 _20156_ (.A1(_03731_),
    .A2(_03759_),
    .ZN(_14790_));
 NOR2_X1 _20157_ (.A1(_03740_),
    .A2(_03753_),
    .ZN(_14792_));
 NOR2_X1 _20158_ (.A1(_03748_),
    .A2(_03745_),
    .ZN(_14791_));
 NAND2_X1 _20159_ (.A1(_03739_),
    .A2(net431),
    .ZN(_14800_));
 NAND2_X1 _20160_ (.A1(net321),
    .A2(_03771_),
    .ZN(_14809_));
 NOR2_X1 _20161_ (.A1(_03692_),
    .A2(_03792_),
    .ZN(_14813_));
 BUF_X2 _20162_ (.A(_00814_),
    .Z(_03808_));
 OAI21_X1 _20163_ (.A(_03803_),
    .B1(_03795_),
    .B2(_03808_),
    .ZN(_03809_));
 AND2_X1 _20164_ (.A1(_03785_),
    .A2(_03809_),
    .ZN(_14824_));
 NAND2_X1 _20165_ (.A1(_03712_),
    .A2(_03781_),
    .ZN(_14842_));
 NOR2_X1 _20166_ (.A1(_03740_),
    .A2(_03759_),
    .ZN(_14849_));
 NOR2_X1 _20167_ (.A1(_03748_),
    .A2(_03753_),
    .ZN(_14848_));
 NOR2_X1 _20168_ (.A1(_03746_),
    .A2(_03754_),
    .ZN(_14847_));
 NAND2_X1 _20169_ (.A1(_03739_),
    .A2(_03756_),
    .ZN(_14856_));
 NAND2_X1 _20170_ (.A1(net321),
    .A2(_03777_),
    .ZN(_14865_));
 NAND2_X2 _20171_ (.A1(_03697_),
    .A2(_03798_),
    .ZN(_14866_));
 INV_X1 _20172_ (.A(_14866_),
    .ZN(_14971_));
 INV_X1 _20173_ (.A(_00845_),
    .ZN(_03810_));
 NAND2_X1 _20174_ (.A1(_03810_),
    .A2(_11434_),
    .ZN(_03811_));
 AOI21_X1 _20175_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03811_),
    .ZN(_14876_));
 NAND2_X1 _20176_ (.A1(_03722_),
    .A2(_03781_),
    .ZN(_14897_));
 NOR2_X1 _20177_ (.A1(_03748_),
    .A2(_03759_),
    .ZN(_14901_));
 NOR2_X1 _20178_ (.A1(_03754_),
    .A2(_03753_),
    .ZN(_14900_));
 NOR2_X1 _20179_ (.A1(_03746_),
    .A2(_03761_),
    .ZN(_14902_));
 NAND2_X1 _20180_ (.A1(_03739_),
    .A2(_03764_),
    .ZN(_14909_));
 BUF_X4 _20181_ (.A(_03784_),
    .Z(_03812_));
 NAND2_X1 _20182_ (.A1(net321),
    .A2(_03812_),
    .ZN(_14919_));
 NAND2_X1 _20183_ (.A1(net324),
    .A2(_03798_),
    .ZN(_14918_));
 INV_X1 _20184_ (.A(_14918_),
    .ZN(_14972_));
 BUF_X2 _20185_ (.A(_00876_),
    .Z(_03813_));
 OAI21_X1 _20186_ (.A(_03803_),
    .B1(_03795_),
    .B2(_03813_),
    .ZN(_03814_));
 AND2_X1 _20187_ (.A1(_03785_),
    .A2(_03814_),
    .ZN(_14931_));
 NAND2_X1 _20188_ (.A1(_03731_),
    .A2(_03781_),
    .ZN(_14950_));
 NAND2_X1 _20189_ (.A1(net431),
    .A2(_03767_),
    .ZN(_14954_));
 NAND2_X1 _20190_ (.A1(_03739_),
    .A2(_03771_),
    .ZN(_14963_));
 AND2_X1 _20191_ (.A1(net322),
    .A2(_03798_),
    .ZN(_14973_));
 BUF_X2 _20192_ (.A(_00907_),
    .Z(_03815_));
 OAI21_X1 _20193_ (.A(_03803_),
    .B1(_03795_),
    .B2(_03815_),
    .ZN(_03816_));
 AND2_X1 _20194_ (.A1(_03785_),
    .A2(_03816_),
    .ZN(_14984_));
 NAND2_X1 _20195_ (.A1(_03740_),
    .A2(net364),
    .ZN(_15002_));
 NAND2_X1 _20196_ (.A1(_03756_),
    .A2(_03767_),
    .ZN(_15009_));
 NAND2_X1 _20197_ (.A1(_03739_),
    .A2(_03777_),
    .ZN(_15015_));
 NAND2_X1 _20198_ (.A1(_03717_),
    .A2(_03798_),
    .ZN(_15016_));
 INV_X1 _20199_ (.A(_15016_),
    .ZN(_15105_));
 BUF_X2 _20200_ (.A(_00938_),
    .Z(_03817_));
 OAI21_X1 _20201_ (.A(_03802_),
    .B1(_03795_),
    .B2(_03817_),
    .ZN(_03818_));
 AND2_X1 _20202_ (.A1(_03785_),
    .A2(_03818_),
    .ZN(_15030_));
 NAND2_X1 _20203_ (.A1(_03748_),
    .A2(_03781_),
    .ZN(_15050_));
 NAND2_X1 _20204_ (.A1(_03767_),
    .A2(_03764_),
    .ZN(_15053_));
 NAND2_X1 _20205_ (.A1(_03739_),
    .A2(_03812_),
    .ZN(_15061_));
 NAND2_X1 _20206_ (.A1(_03729_),
    .A2(_03798_),
    .ZN(_15060_));
 INV_X1 _20207_ (.A(_15060_),
    .ZN(_15103_));
 BUF_X2 _20208_ (.A(_00969_),
    .Z(_03819_));
 OAI21_X1 _20209_ (.A(_03802_),
    .B1(_03795_),
    .B2(_03819_),
    .ZN(_03820_));
 AND2_X1 _20210_ (.A1(_03785_),
    .A2(_03820_),
    .ZN(_15073_));
 NAND2_X1 _20211_ (.A1(_03754_),
    .A2(net364),
    .ZN(_15093_));
 NAND2_X1 _20212_ (.A1(_03767_),
    .A2(_03771_),
    .ZN(_15098_));
 AND2_X1 _20213_ (.A1(_03738_),
    .A2(_03798_),
    .ZN(_15104_));
 INV_X1 _20214_ (.A(_01000_),
    .ZN(_03821_));
 NAND2_X1 _20215_ (.A1(_03821_),
    .A2(_11434_),
    .ZN(_03822_));
 AOI21_X2 _20216_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03822_),
    .ZN(_15117_));
 NAND2_X1 _20217_ (.A1(_03761_),
    .A2(net364),
    .ZN(_15136_));
 NAND2_X1 _20218_ (.A1(_03767_),
    .A2(_03777_),
    .ZN(_15141_));
 INV_X2 _20219_ (.A(_03745_),
    .ZN(_03823_));
 NAND2_X1 _20220_ (.A1(_03823_),
    .A2(_03798_),
    .ZN(_15142_));
 INV_X1 _20221_ (.A(_15142_),
    .ZN(_15218_));
 CLKBUF_X3 _20222_ (.A(_01031_),
    .Z(_03824_));
 OAI21_X1 _20223_ (.A(_03802_),
    .B1(_03795_),
    .B2(_03824_),
    .ZN(_03825_));
 AND2_X1 _20224_ (.A1(_03785_),
    .A2(_03825_),
    .ZN(_15156_));
 NAND2_X1 _20225_ (.A1(_03768_),
    .A2(net364),
    .ZN(_15175_));
 NAND2_X1 _20226_ (.A1(_03767_),
    .A2(_03812_),
    .ZN(_15179_));
 INV_X2 _20227_ (.A(_03752_),
    .ZN(_03826_));
 NAND2_X1 _20228_ (.A1(_03826_),
    .A2(_03797_),
    .ZN(_15180_));
 INV_X1 _20229_ (.A(_15180_),
    .ZN(_15217_));
 BUF_X2 _20230_ (.A(_01062_),
    .Z(_03827_));
 OAI21_X1 _20231_ (.A(_03802_),
    .B1(_03795_),
    .B2(_03827_),
    .ZN(_03828_));
 AND2_X1 _20232_ (.A1(_03785_),
    .A2(_03828_),
    .ZN(_15193_));
 NAND2_X1 _20233_ (.A1(_03775_),
    .A2(net335),
    .ZN(_15212_));
 NOR2_X1 _20234_ (.A1(_03759_),
    .A2(_03792_),
    .ZN(_15216_));
 INV_X1 _20235_ (.A(_01093_),
    .ZN(_03829_));
 NAND2_X1 _20236_ (.A1(_03829_),
    .A2(_11434_),
    .ZN(_03830_));
 AOI21_X1 _20237_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03830_),
    .ZN(_15232_));
 NAND2_X1 _20238_ (.A1(_03782_),
    .A2(net364),
    .ZN(_15250_));
 INV_X1 _20239_ (.A(_01124_),
    .ZN(_03831_));
 NAND2_X1 _20240_ (.A1(_03831_),
    .A2(_11434_),
    .ZN(_03832_));
 AOI21_X2 _20241_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03832_),
    .ZN(_15272_));
 NAND2_X1 _20242_ (.A1(net364),
    .A2(_03796_),
    .ZN(_15290_));
 OAI21_X1 _20243_ (.A(_03802_),
    .B1(_03794_),
    .B2(_03412_),
    .ZN(_03833_));
 AND2_X1 _20244_ (.A1(_03785_),
    .A2(_03833_),
    .ZN(_15308_));
 NAND2_X1 _20245_ (.A1(net364),
    .A2(_03792_),
    .ZN(_15325_));
 NAND2_X1 _20246_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(_11434_),
    .ZN(_03834_));
 AOI21_X2 _20247_ (.A(_03720_),
    .B1(_03803_),
    .B2(_03834_),
    .ZN(_15337_));
 INV_X1 _20248_ (.A(_15327_),
    .ZN(_15328_));
 INV_X1 _20249_ (.A(_15220_),
    .ZN(_15221_));
 INV_X4 _20250_ (.A(_14815_),
    .ZN(_14880_));
 NAND4_X2 _20251_ (.A1(_10304_),
    .A2(_10522_),
    .A3(_10670_),
    .A4(_10997_),
    .ZN(_03835_));
 OR4_X2 _20252_ (.A1(_03465_),
    .A2(_10886_),
    .A3(_10876_),
    .A4(_03835_),
    .ZN(_03836_));
 OR2_X2 _20253_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.load_err_q ),
    .ZN(_03837_));
 NOR2_X4 _20254_ (.A1(\id_stage_i.controller_i.exc_req_q ),
    .A2(_03837_),
    .ZN(_03838_));
 OR4_X2 _20255_ (.A1(_10886_),
    .A2(_10887_),
    .A3(_10889_),
    .A4(_03835_),
    .ZN(_03839_));
 OAI211_X2 _20256_ (.A(_03836_),
    .B(_03838_),
    .C1(_03465_),
    .C2(_03839_),
    .ZN(_03840_));
 OR3_X1 _20257_ (.A1(_03465_),
    .A2(_10892_),
    .A3(_10876_),
    .ZN(_03841_));
 BUF_X2 _20258_ (.A(_01157_),
    .Z(_03842_));
 NAND2_X2 _20259_ (.A1(_10304_),
    .A2(_11419_),
    .ZN(_03843_));
 BUF_X4 _20260_ (.A(_01156_),
    .Z(_03844_));
 NAND2_X1 _20261_ (.A1(_03462_),
    .A2(_03463_),
    .ZN(_03845_));
 INV_X1 _20262_ (.A(\cs_registers_i.dcsr_q[15] ),
    .ZN(_03846_));
 OR2_X1 _20263_ (.A1(_03462_),
    .A2(_03463_),
    .ZN(_03847_));
 INV_X1 _20264_ (.A(\cs_registers_i.dcsr_q[12] ),
    .ZN(_03848_));
 OAI221_X2 _20265_ (.A(_03844_),
    .B1(_03845_),
    .B2(_03846_),
    .C1(_03847_),
    .C2(_03848_),
    .ZN(_03849_));
 NAND3_X1 _20266_ (.A1(_03842_),
    .A2(_03843_),
    .A3(_03849_),
    .ZN(_03850_));
 NOR2_X1 _20267_ (.A1(_11419_),
    .A2(\id_stage_i.controller_i.illegal_insn_q ),
    .ZN(_03851_));
 NAND2_X1 _20268_ (.A1(_10466_),
    .A2(_03851_),
    .ZN(_03852_));
 OR2_X1 _20269_ (.A1(_03835_),
    .A2(_03852_),
    .ZN(_03853_));
 OR4_X2 _20270_ (.A1(_03841_),
    .A2(_03838_),
    .A3(_03850_),
    .A4(_03853_),
    .ZN(_03854_));
 NAND3_X2 _20271_ (.A1(_03461_),
    .A2(_03840_),
    .A3(_03854_),
    .ZN(_03855_));
 AOI22_X4 _20272_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net145),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net146),
    .ZN(_03856_));
 AOI22_X4 _20273_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net147),
    .B1(\cs_registers_i.mie_q[7] ),
    .B2(net148),
    .ZN(_03857_));
 AOI22_X4 _20274_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net143),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net144),
    .ZN(_03858_));
 AOI22_X4 _20275_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net136),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net142),
    .ZN(_03859_));
 AND4_X1 _20276_ (.A1(_03856_),
    .A2(_03857_),
    .A3(_03858_),
    .A4(_03859_),
    .ZN(_03860_));
 AOI22_X2 _20277_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net137),
    .B1(\cs_registers_i.mie_q[11] ),
    .B2(net138),
    .ZN(_03861_));
 AOI22_X2 _20278_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net149),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net150),
    .ZN(_03862_));
 AOI22_X4 _20279_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net139),
    .B1(\cs_registers_i.mie_q[13] ),
    .B2(net140),
    .ZN(_03863_));
 NAND2_X2 _20280_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(net141),
    .ZN(_03864_));
 AND4_X1 _20281_ (.A1(_03861_),
    .A2(_03862_),
    .A3(_03863_),
    .A4(_03864_),
    .ZN(_03865_));
 AOI22_X4 _20282_ (.A1(net135),
    .A2(\cs_registers_i.mie_q[15] ),
    .B1(\cs_registers_i.mie_q[17] ),
    .B2(net151),
    .ZN(_03866_));
 BUF_X2 _20283_ (.A(irq_nm_i),
    .Z(_03867_));
 AOI21_X2 _20284_ (.A(_03867_),
    .B1(\cs_registers_i.mie_q[16] ),
    .B2(net152),
    .ZN(_03868_));
 NAND4_X4 _20285_ (.A1(_03860_),
    .A2(_03865_),
    .A3(_03866_),
    .A4(_03868_),
    .ZN(_03869_));
 BUF_X4 _20286_ (.A(\cs_registers_i.nmi_mode_i ),
    .Z(_03870_));
 NOR2_X1 _20287_ (.A1(_03867_),
    .A2(\cs_registers_i.csr_mstatus_mie_o ),
    .ZN(_03871_));
 NOR3_X4 _20288_ (.A1(_03477_),
    .A2(_03870_),
    .A3(_03871_),
    .ZN(_03872_));
 NAND4_X4 _20289_ (.A1(_11420_),
    .A2(_03459_),
    .A3(_03869_),
    .A4(_03872_),
    .ZN(_03873_));
 NAND3_X1 _20290_ (.A1(\id_stage_i.branch_set ),
    .A2(net22),
    .A3(_03843_),
    .ZN(_03874_));
 INV_X2 _20291_ (.A(_11422_),
    .ZN(_03875_));
 NAND3_X4 _20292_ (.A1(_03458_),
    .A2(_03875_),
    .A3(_11424_),
    .ZN(_03876_));
 NAND2_X4 _20293_ (.A1(_03458_),
    .A2(_11424_),
    .ZN(_03877_));
 NOR2_X4 _20294_ (.A1(_03875_),
    .A2(_03877_),
    .ZN(_03878_));
 CLKBUF_X2 _20295_ (.A(\cs_registers_i.dcsr_q[2] ),
    .Z(_03879_));
 OR2_X2 _20296_ (.A1(_03879_),
    .A2(net69),
    .ZN(_03880_));
 OAI21_X2 _20297_ (.A(_03878_),
    .B1(_03880_),
    .B2(_11420_),
    .ZN(_03881_));
 AND4_X2 _20298_ (.A1(_03873_),
    .A2(_03874_),
    .A3(_03876_),
    .A4(_03881_),
    .ZN(_03882_));
 NAND2_X2 _20299_ (.A1(_03855_),
    .A2(_03882_),
    .ZN(_03883_));
 AOI21_X2 _20300_ (.A(_10352_),
    .B1(_10342_),
    .B2(_10349_),
    .ZN(_03884_));
 NOR2_X2 _20301_ (.A1(_10340_),
    .A2(_03884_),
    .ZN(_03885_));
 NOR3_X4 _20302_ (.A1(_10306_),
    .A2(_10401_),
    .A3(_03438_),
    .ZN(_03886_));
 NAND4_X4 _20303_ (.A1(net22),
    .A2(_03843_),
    .A3(_03885_),
    .A4(_03886_),
    .ZN(_03887_));
 NOR2_X2 _20304_ (.A1(_03434_),
    .A2(_03887_),
    .ZN(_03888_));
 NOR2_X2 _20305_ (.A1(_03883_),
    .A2(_03888_),
    .ZN(_03889_));
 NAND3_X4 _20306_ (.A1(_03458_),
    .A2(_11422_),
    .A3(_11424_),
    .ZN(_03890_));
 OR2_X2 _20307_ (.A1(\id_stage_i.controller_i.exc_req_q ),
    .A2(_03837_),
    .ZN(_03891_));
 OAI21_X2 _20308_ (.A(_03459_),
    .B1(_03891_),
    .B2(_11420_),
    .ZN(_03892_));
 NAND2_X4 _20309_ (.A1(_03890_),
    .A2(_03892_),
    .ZN(_03893_));
 NAND2_X4 _20310_ (.A1(_03466_),
    .A2(_03468_),
    .ZN(_03894_));
 NAND3_X4 _20311_ (.A1(_10661_),
    .A2(_03475_),
    .A3(_03468_),
    .ZN(_03895_));
 OAI21_X2 _20312_ (.A(_03894_),
    .B1(_03895_),
    .B2(_03891_),
    .ZN(_03896_));
 AOI221_X2 _20313_ (.A(_03893_),
    .B1(_03896_),
    .B2(_03461_),
    .C1(_11425_),
    .C2(_11420_),
    .ZN(_03897_));
 NOR2_X1 _20314_ (.A1(_03889_),
    .A2(_03897_),
    .ZN(_03898_));
 NAND4_X4 _20315_ (.A1(_03856_),
    .A2(_03857_),
    .A3(_03858_),
    .A4(_03859_),
    .ZN(_03899_));
 AND2_X1 _20316_ (.A1(_03861_),
    .A2(_03862_),
    .ZN(_03900_));
 NAND3_X2 _20317_ (.A1(_03900_),
    .A2(_03863_),
    .A3(_03864_),
    .ZN(_03901_));
 NOR2_X4 _20318_ (.A1(_03899_),
    .A2(_03901_),
    .ZN(_03902_));
 NAND2_X1 _20319_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(net140),
    .ZN(_03903_));
 AND2_X1 _20320_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net139),
    .ZN(_03904_));
 NAND2_X1 _20321_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net148),
    .ZN(_03905_));
 NAND2_X1 _20322_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net147),
    .ZN(_03906_));
 NAND2_X1 _20323_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(net144),
    .ZN(_03907_));
 NAND2_X1 _20324_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net143),
    .ZN(_03908_));
 NAND3_X1 _20325_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net142),
    .A3(_03908_),
    .ZN(_03909_));
 AOI22_X1 _20326_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net145),
    .B1(_03907_),
    .B2(_03909_),
    .ZN(_03910_));
 AND2_X1 _20327_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net146),
    .ZN(_03911_));
 OAI21_X1 _20328_ (.A(_03906_),
    .B1(_03910_),
    .B2(_03911_),
    .ZN(_03912_));
 AOI22_X1 _20329_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net149),
    .B1(_03905_),
    .B2(_03912_),
    .ZN(_03913_));
 AOI21_X1 _20330_ (.A(_03913_),
    .B1(net150),
    .B2(\cs_registers_i.mie_q[9] ),
    .ZN(_03914_));
 AOI21_X1 _20331_ (.A(_03914_),
    .B1(net137),
    .B2(\cs_registers_i.mie_q[10] ),
    .ZN(_03915_));
 AOI21_X1 _20332_ (.A(_03915_),
    .B1(net138),
    .B2(\cs_registers_i.mie_q[11] ),
    .ZN(_03916_));
 OAI21_X1 _20333_ (.A(_03903_),
    .B1(_03904_),
    .B2(_03916_),
    .ZN(_03917_));
 INV_X2 _20334_ (.A(_03870_),
    .ZN(_03918_));
 AOI221_X2 _20335_ (.A(_03902_),
    .B1(_03917_),
    .B2(_03864_),
    .C1(_03867_),
    .C2(_03918_),
    .ZN(_03919_));
 NOR2_X2 _20336_ (.A1(_03873_),
    .A2(_03919_),
    .ZN(_03920_));
 NAND2_X4 _20337_ (.A1(_03461_),
    .A2(_03838_),
    .ZN(_03921_));
 NOR2_X4 _20338_ (.A1(_03894_),
    .A2(_03921_),
    .ZN(_03922_));
 BUF_X4 _20339_ (.A(_03922_),
    .Z(_03923_));
 BUF_X4 _20340_ (.A(_03923_),
    .Z(_03924_));
 NOR2_X4 _20341_ (.A1(_03895_),
    .A2(_03921_),
    .ZN(_03925_));
 BUF_X4 _20342_ (.A(_03925_),
    .Z(_03926_));
 BUF_X4 _20343_ (.A(_03926_),
    .Z(_03927_));
 AOI221_X2 _20344_ (.A(_03920_),
    .B1(_03924_),
    .B2(\cs_registers_i.csr_mepc_o[2] ),
    .C1(_03927_),
    .C2(\cs_registers_i.csr_depc_o[2] ),
    .ZN(_03928_));
 BUF_X4 _20345_ (.A(net22),
    .Z(_03929_));
 BUF_X4 _20346_ (.A(_03929_),
    .Z(_03930_));
 BUF_X4 _20347_ (.A(_03930_),
    .Z(_03931_));
 NAND2_X1 _20348_ (.A1(_03931_),
    .A2(\alu_adder_result_ex[2] ),
    .ZN(_03932_));
 NAND2_X1 _20349_ (.A1(_03928_),
    .A2(_03932_),
    .ZN(_03933_));
 NAND2_X2 _20350_ (.A1(_03898_),
    .A2(_03933_),
    .ZN(_03934_));
 OAI211_X4 _20351_ (.A(_03855_),
    .B(_03882_),
    .C1(_03887_),
    .C2(_03434_),
    .ZN(_03935_));
 BUF_X4 _20352_ (.A(_03935_),
    .Z(_03936_));
 CLKBUF_X3 _20353_ (.A(_03936_),
    .Z(_03937_));
 BUF_X4 _20354_ (.A(_03937_),
    .Z(_03938_));
 BUF_X4 _20355_ (.A(_03938_),
    .Z(_03939_));
 INV_X1 _20356_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .ZN(_03940_));
 OAI21_X2 _20357_ (.A(_03934_),
    .B1(_03939_),
    .B2(_03940_),
    .ZN(_16108_));
 INV_X1 _20358_ (.A(_03873_),
    .ZN(_03941_));
 INV_X1 _20359_ (.A(_03863_),
    .ZN(_03942_));
 INV_X1 _20360_ (.A(_03856_),
    .ZN(_03943_));
 OAI21_X1 _20361_ (.A(_03857_),
    .B1(_03858_),
    .B2(_03943_),
    .ZN(_03944_));
 NAND2_X1 _20362_ (.A1(_03862_),
    .A2(_03944_),
    .ZN(_03945_));
 AOI21_X1 _20363_ (.A(_03942_),
    .B1(_03945_),
    .B2(_03861_),
    .ZN(_03946_));
 INV_X1 _20364_ (.A(_03867_),
    .ZN(_03947_));
 OAI221_X2 _20365_ (.A(_03864_),
    .B1(_03901_),
    .B2(_03899_),
    .C1(_03947_),
    .C2(_03870_),
    .ZN(_03948_));
 OAI21_X2 _20366_ (.A(_03941_),
    .B1(_03946_),
    .B2(_03948_),
    .ZN(_03949_));
 INV_X1 _20367_ (.A(_01163_),
    .ZN(_03950_));
 AOI22_X1 _20368_ (.A1(net22),
    .A2(\alu_adder_result_ex[3] ),
    .B1(_03925_),
    .B2(_03950_),
    .ZN(_03951_));
 NAND2_X2 _20369_ (.A1(_03436_),
    .A2(_03459_),
    .ZN(_03952_));
 NOR2_X4 _20370_ (.A1(_03952_),
    .A2(_03838_),
    .ZN(_03953_));
 INV_X2 _20371_ (.A(_03844_),
    .ZN(_03954_));
 AOI22_X1 _20372_ (.A1(\cs_registers_i.csr_mepc_o[3] ),
    .A2(_03922_),
    .B1(_03953_),
    .B2(_03954_),
    .ZN(_03955_));
 AND4_X2 _20373_ (.A1(_03935_),
    .A2(_03949_),
    .A3(_03951_),
    .A4(_03955_),
    .ZN(_03956_));
 BUF_X4 _20374_ (.A(_03889_),
    .Z(_03957_));
 INV_X1 _20375_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .ZN(_03958_));
 AOI21_X2 _20376_ (.A(_03956_),
    .B1(_03957_),
    .B2(_03958_),
    .ZN(_16110_));
 BUF_X4 _20377_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Z(_03959_));
 OAI21_X1 _20378_ (.A(_03959_),
    .B1(_03939_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .ZN(_03960_));
 INV_X1 _20379_ (.A(_03960_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 BUF_X4 _20380_ (.A(\cs_registers_i.pc_if_i[1] ),
    .Z(_03961_));
 CLKBUF_X3 _20381_ (.A(_03961_),
    .Z(_03962_));
 BUF_X4 _20382_ (.A(_03962_),
    .Z(_03963_));
 BUF_X2 _20383_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_03964_));
 INV_X4 _20384_ (.A(_03964_),
    .ZN(_03965_));
 BUF_X2 _20385_ (.A(instr_err_i),
    .Z(_03966_));
 CLKBUF_X2 _20386_ (.A(instr_rdata_i[17]),
    .Z(_03967_));
 CLKBUF_X2 _20387_ (.A(instr_rdata_i[16]),
    .Z(_03968_));
 AOI21_X1 _20388_ (.A(_03966_),
    .B1(_03967_),
    .B2(_03968_),
    .ZN(_03969_));
 AND2_X1 _20389_ (.A1(_03965_),
    .A2(_03969_),
    .ZN(_03970_));
 BUF_X2 _20390_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .Z(_03971_));
 AOI21_X2 _20391_ (.A(_03971_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .ZN(_03972_));
 BUF_X4 _20392_ (.A(_03964_),
    .Z(_03973_));
 AOI21_X4 _20393_ (.A(_03970_),
    .B1(_03972_),
    .B2(_03973_),
    .ZN(_03974_));
 NAND2_X2 _20394_ (.A1(_03963_),
    .A2(_03974_),
    .ZN(_03975_));
 AOI21_X1 _20395_ (.A(_03966_),
    .B1(net113),
    .B2(net104),
    .ZN(_03976_));
 AOI21_X1 _20396_ (.A(_03971_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .ZN(_03977_));
 BUF_X4 _20397_ (.A(_03973_),
    .Z(_03978_));
 CLKBUF_X3 _20398_ (.A(_03978_),
    .Z(_03979_));
 MUX2_X2 _20399_ (.A(_03976_),
    .B(_03977_),
    .S(_03979_),
    .Z(_03980_));
 BUF_X4 _20400_ (.A(_03963_),
    .Z(_03981_));
 OAI21_X4 _20401_ (.A(_03975_),
    .B1(_03980_),
    .B2(_03981_),
    .ZN(_15831_));
 INV_X1 _20402_ (.A(_15831_),
    .ZN(_15353_));
 INV_X1 _20403_ (.A(net154),
    .ZN(_03982_));
 OR2_X1 _20404_ (.A1(net69),
    .A2(core_busy_q),
    .ZN(_03983_));
 OAI21_X2 _20405_ (.A(fetch_enable_q),
    .B1(_03869_),
    .B2(_03983_),
    .ZN(net155));
 AND2_X1 _20406_ (.A1(_03982_),
    .A2(net155),
    .ZN(_03984_));
 INV_X1 _20407_ (.A(_03984_),
    .ZN(_00006_));
 BUF_X8 _20408_ (.A(_03661_),
    .Z(_03985_));
 NAND2_X1 _20409_ (.A1(net354),
    .A2(_03689_),
    .ZN(_14074_));
 BUF_X4 _20410_ (.A(_03658_),
    .Z(_03986_));
 NOR2_X1 _20411_ (.A1(_03806_),
    .A2(_03669_),
    .ZN(_03987_));
 CLKBUF_X3 _20412_ (.A(_11433_),
    .Z(_03988_));
 AOI21_X1 _20413_ (.A(_03987_),
    .B1(_03988_),
    .B2(_00557_),
    .ZN(_03989_));
 BUF_X4 _20414_ (.A(_11431_),
    .Z(_03990_));
 AOI22_X2 _20415_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_03986_),
    .B1(_03989_),
    .B2(_03990_),
    .ZN(_14079_));
 NAND2_X1 _20416_ (.A1(_03985_),
    .A2(_03702_),
    .ZN(_14089_));
 INV_X1 _20417_ (.A(_15577_),
    .ZN(_14099_));
 NOR2_X1 _20418_ (.A1(_03810_),
    .A2(_03669_),
    .ZN(_03991_));
 AOI21_X1 _20419_ (.A(_03991_),
    .B1(_03988_),
    .B2(_00559_),
    .ZN(_03992_));
 AOI22_X2 _20420_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_03986_),
    .B1(_03992_),
    .B2(_03990_),
    .ZN(_14109_));
 INV_X1 _20421_ (.A(_15585_),
    .ZN(_14117_));
 NAND2_X1 _20422_ (.A1(_03683_),
    .A2(net324),
    .ZN(_14145_));
 NAND2_X1 _20423_ (.A1(_03985_),
    .A2(_03726_),
    .ZN(_14159_));
 INV_X1 _20424_ (.A(_15614_),
    .ZN(_14172_));
 NAND2_X1 _20425_ (.A1(_03690_),
    .A2(_03703_),
    .ZN(_14177_));
 INV_X1 _20426_ (.A(_15633_),
    .ZN(_14229_));
 INV_X1 _20427_ (.A(_15651_),
    .ZN(_14269_));
 INV_X1 _20428_ (.A(_15664_),
    .ZN(_14312_));
 BUF_X8 _20429_ (.A(_03729_),
    .Z(_03993_));
 NAND2_X1 _20430_ (.A1(_03695_),
    .A2(_03993_),
    .ZN(_14326_));
 NAND2_X1 _20431_ (.A1(net354),
    .A2(_03764_),
    .ZN(_14352_));
 BUF_X8 _20432_ (.A(_03703_),
    .Z(_03994_));
 NAND2_X1 _20433_ (.A1(_03994_),
    .A2(_03726_),
    .ZN(_14385_));
 NAND2_X1 _20434_ (.A1(_03695_),
    .A2(_03823_),
    .ZN(_14428_));
 NAND2_X1 _20435_ (.A1(_03708_),
    .A2(_03993_),
    .ZN(_14433_));
 NAND2_X1 _20436_ (.A1(_03994_),
    .A2(_03735_),
    .ZN(_14441_));
 BUF_X8 _20437_ (.A(_03717_),
    .Z(_03995_));
 NAND2_X1 _20438_ (.A1(_03995_),
    .A2(_03726_),
    .ZN(_14487_));
 NAND2_X2 _20439_ (.A1(_03994_),
    .A2(_03742_),
    .ZN(_14499_));
 NAND2_X1 _20440_ (.A1(net354),
    .A2(_03812_),
    .ZN(_14518_));
 NAND2_X1 _20441_ (.A1(_03726_),
    .A2(_03729_),
    .ZN(_14553_));
 BUF_X4 _20442_ (.A(_03774_),
    .Z(_03996_));
 NAND2_X1 _20443_ (.A1(_03690_),
    .A2(_03996_),
    .ZN(_14609_));
 NAND2_X1 _20444_ (.A1(_03995_),
    .A2(_03742_),
    .ZN(_14622_));
 NAND2_X1 _20445_ (.A1(net323),
    .A2(_03756_),
    .ZN(_14633_));
 NOR2_X2 clone2 (.A1(_03792_),
    .A2(_03662_),
    .ZN(net2));
 NAND2_X1 _20447_ (.A1(_03702_),
    .A2(_03765_),
    .ZN(_14669_));
 NAND2_X1 _20448_ (.A1(_03993_),
    .A2(_03742_),
    .ZN(_14682_));
 BUF_X8 _20449_ (.A(_03697_),
    .Z(_03998_));
 NAND2_X1 _20450_ (.A1(net325),
    .A2(_03771_),
    .ZN(_14692_));
 NAND2_X1 _20451_ (.A1(_03708_),
    .A2(_03765_),
    .ZN(_14727_));
 NAND2_X1 _20452_ (.A1(_03993_),
    .A2(net431),
    .ZN(_14740_));
 NAND2_X1 _20453_ (.A1(net325),
    .A2(_03777_),
    .ZN(_14750_));
 NAND2_X1 _20454_ (.A1(_03708_),
    .A2(_03996_),
    .ZN(_14785_));
 NAND2_X1 _20455_ (.A1(net337),
    .A2(_03764_),
    .ZN(_14798_));
 NAND2_X1 _20456_ (.A1(net323),
    .A2(_03777_),
    .ZN(_14808_));
 NAND2_X1 _20457_ (.A1(_03993_),
    .A2(_03764_),
    .ZN(_14855_));
 NAND2_X1 _20458_ (.A1(_03735_),
    .A2(net291),
    .ZN(_14895_));
 NAND2_X1 _20459_ (.A1(_03993_),
    .A2(_03771_),
    .ZN(_14908_));
 NAND2_X1 _20460_ (.A1(_03735_),
    .A2(_03996_),
    .ZN(_14949_));
 NAND2_X1 _20461_ (.A1(net337),
    .A2(_03812_),
    .ZN(_14961_));
 NAND2_X1 _20462_ (.A1(_03823_),
    .A2(_03771_),
    .ZN(_15007_));
 NAND2_X1 _20463_ (.A1(_03993_),
    .A2(_03812_),
    .ZN(_15014_));
 INV_X1 _20464_ (.A(_14975_),
    .ZN(_14976_));
 NAND2_X1 _20465_ (.A1(_03756_),
    .A2(net291),
    .ZN(_15048_));
 NAND2_X1 _20466_ (.A1(_03764_),
    .A2(net291),
    .ZN(_15091_));
 NAND2_X1 _20467_ (.A1(_03823_),
    .A2(_03812_),
    .ZN(_15096_));
 NAND2_X1 _20468_ (.A1(_03764_),
    .A2(_03996_),
    .ZN(_15135_));
 NAND2_X1 _20469_ (.A1(_03826_),
    .A2(_03812_),
    .ZN(_15140_));
 NAND2_X1 _20470_ (.A1(_03771_),
    .A2(_03996_),
    .ZN(_15174_));
 NAND2_X1 _20471_ (.A1(_03996_),
    .A2(_03777_),
    .ZN(_15211_));
 INV_X4 _20472_ (.A(_15024_),
    .ZN(_15025_));
 NAND2_X2 _20473_ (.A1(net291),
    .A2(_03798_),
    .ZN(_15251_));
 NAND2_X1 _20474_ (.A1(net354),
    .A2(_03683_),
    .ZN(_14070_));
 CLKBUF_X2 _20475_ (.A(_11402_),
    .Z(_03999_));
 OR2_X1 _20476_ (.A1(_00556_),
    .A2(_03999_),
    .ZN(_04000_));
 OAI21_X1 _20477_ (.A(_04000_),
    .B1(_03988_),
    .B2(_03804_),
    .ZN(_04001_));
 AOI22_X2 _20478_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_03986_),
    .B1(_04001_),
    .B2(_03990_),
    .ZN(_14075_));
 OR2_X1 _20479_ (.A1(_00558_),
    .A2(_03999_),
    .ZN(_04002_));
 OAI21_X1 _20480_ (.A(_04002_),
    .B1(_03988_),
    .B2(_03808_),
    .ZN(_04003_));
 AOI22_X2 _20481_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_03986_),
    .B1(_04003_),
    .B2(_03990_),
    .ZN(_14090_));
 NAND2_X1 _20482_ (.A1(net354),
    .A2(_03715_),
    .ZN(_14133_));
 INV_X1 _20483_ (.A(_15595_),
    .ZN(_14141_));
 OR2_X1 _20484_ (.A1(_00561_),
    .A2(_03999_),
    .ZN(_04004_));
 OAI21_X1 _20485_ (.A(_04004_),
    .B1(_03988_),
    .B2(_03815_),
    .ZN(_04005_));
 AOI22_X2 _20486_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_03986_),
    .B1(_04005_),
    .B2(_03990_),
    .ZN(_14160_));
 INV_X1 _20487_ (.A(_15606_),
    .ZN(_14168_));
 NAND2_X1 _20488_ (.A1(_03985_),
    .A2(_03735_),
    .ZN(_14191_));
 INV_X1 _20489_ (.A(_15620_),
    .ZN(_14199_));
 NAND2_X1 _20490_ (.A1(_03998_),
    .A2(_03702_),
    .ZN(_14209_));
 NAND2_X1 _20491_ (.A1(_03985_),
    .A2(_03742_),
    .ZN(_14222_));
 INV_X1 _20492_ (.A(_15639_),
    .ZN(_14230_));
 NAND2_X1 _20493_ (.A1(_03690_),
    .A2(_03995_),
    .ZN(_14244_));
 NAND2_X1 _20494_ (.A1(_03998_),
    .A2(_03708_),
    .ZN(_14249_));
 NAND2_X1 _20495_ (.A1(_03985_),
    .A2(_03749_),
    .ZN(_14262_));
 INV_X1 _20496_ (.A(_15655_),
    .ZN(_14270_));
 NAND2_X1 _20497_ (.A1(_03695_),
    .A2(net336),
    .ZN(_14284_));
 NAND2_X1 _20498_ (.A1(_03998_),
    .A2(_03715_),
    .ZN(_14289_));
 NAND2_X1 _20499_ (.A1(_03661_),
    .A2(_03756_),
    .ZN(_14305_));
 INV_X1 _20500_ (.A(_15668_),
    .ZN(_14313_));
 NAND2_X1 _20501_ (.A1(_03998_),
    .A2(_03726_),
    .ZN(_14332_));
 OR2_X1 _20502_ (.A1(_00566_),
    .A2(_03999_),
    .ZN(_04006_));
 OAI21_X2 _20503_ (.A(_04006_),
    .B1(_03988_),
    .B2(_03827_),
    .ZN(_04007_));
 AOI22_X4 _20504_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(_03986_),
    .B1(_04007_),
    .B2(_03990_),
    .ZN(_14353_));
 NAND2_X1 _20505_ (.A1(_03708_),
    .A2(net336),
    .ZN(_14378_));
 NAND2_X1 _20506_ (.A1(_03661_),
    .A2(_03771_),
    .ZN(_14407_));
 NAND2_X1 _20507_ (.A1(_03690_),
    .A2(_03826_),
    .ZN(_14429_));
 NAND2_X1 _20508_ (.A1(_03661_),
    .A2(_03777_),
    .ZN(_14462_));
 NAND2_X1 _20509_ (.A1(_03715_),
    .A2(_03729_),
    .ZN(_14488_));
 OR2_X1 _20510_ (.A1(_00659_),
    .A2(_03999_),
    .ZN(_04008_));
 OAI21_X1 _20511_ (.A(_04008_),
    .B1(_03988_),
    .B2(_03412_),
    .ZN(_04009_));
 AOI22_X2 _20512_ (.A1(_03408_),
    .A2(_03986_),
    .B1(_04009_),
    .B2(_03990_),
    .ZN(_14519_));
 NAND2_X1 _20513_ (.A1(_03690_),
    .A2(_03765_),
    .ZN(_14540_));
 NAND2_X1 _20514_ (.A1(net325),
    .A2(_03756_),
    .ZN(_14566_));
 NAND2_X1 _20515_ (.A1(_03993_),
    .A2(_03735_),
    .ZN(_14623_));
 NAND2_X1 _20516_ (.A1(_03695_),
    .A2(_03996_),
    .ZN(_14670_));
 NAND2_X1 _20517_ (.A1(net323),
    .A2(_03764_),
    .ZN(_14693_));
 NAND2_X1 _20518_ (.A1(_03702_),
    .A2(_03996_),
    .ZN(_14728_));
 NAND2_X1 _20519_ (.A1(net323),
    .A2(_03771_),
    .ZN(_14751_));
 NAND2_X1 _20520_ (.A1(_03993_),
    .A2(_03756_),
    .ZN(_14799_));
 NAND2_X1 _20521_ (.A1(_03726_),
    .A2(_03765_),
    .ZN(_14843_));
 NAND2_X1 _20522_ (.A1(_03726_),
    .A2(_03774_),
    .ZN(_14896_));
 NAND2_X1 _20523_ (.A1(_03823_),
    .A2(_03763_),
    .ZN(_14955_));
 NAND2_X1 _20524_ (.A1(_03993_),
    .A2(_03777_),
    .ZN(_14962_));
 NAND2_X1 _20525_ (.A1(net431),
    .A2(net291),
    .ZN(_15003_));
 NAND2_X1 _20526_ (.A1(_03826_),
    .A2(_03763_),
    .ZN(_15008_));
 NAND2_X1 _20527_ (.A1(net431),
    .A2(_03774_),
    .ZN(_15049_));
 NAND2_X1 _20528_ (.A1(_03823_),
    .A2(_03777_),
    .ZN(_15054_));
 NAND2_X1 _20529_ (.A1(_03756_),
    .A2(_03774_),
    .ZN(_15092_));
 NAND2_X1 _20530_ (.A1(_03826_),
    .A2(_03776_),
    .ZN(_15097_));
 OR2_X1 _20531_ (.A1(_00185_),
    .A2(_03999_),
    .ZN(_04010_));
 OAI21_X1 _20532_ (.A(_04010_),
    .B1(_03669_),
    .B2(_03800_),
    .ZN(_04011_));
 AOI22_X1 _20533_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A2(_03986_),
    .B1(_04011_),
    .B2(_03990_),
    .ZN(_14071_));
 NAND2_X1 _20534_ (.A1(_03661_),
    .A2(_03694_),
    .ZN(_14081_));
 INV_X1 _20535_ (.A(_15575_),
    .ZN(_14101_));
 NAND2_X1 _20536_ (.A1(_03661_),
    .A2(_03708_),
    .ZN(_14111_));
 INV_X1 _20537_ (.A(_15583_),
    .ZN(_14119_));
 OR2_X1 _20538_ (.A1(_00560_),
    .A2(_03999_),
    .ZN(_04012_));
 OAI21_X1 _20539_ (.A(_04012_),
    .B1(_03669_),
    .B2(_03813_),
    .ZN(_04013_));
 AOI22_X2 _20540_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_03986_),
    .B1(_04013_),
    .B2(_03990_),
    .ZN(_14134_));
 INV_X1 _20541_ (.A(_15597_),
    .ZN(_14142_));
 NAND2_X1 _20542_ (.A1(_03690_),
    .A2(_03697_),
    .ZN(_14147_));
 INV_X1 _20543_ (.A(_15610_),
    .ZN(_14169_));
 INV_X1 _20544_ (.A(_15612_),
    .ZN(_14174_));
 NAND2_X1 _20545_ (.A1(_03695_),
    .A2(_03697_),
    .ZN(_14179_));
 OR2_X1 _20546_ (.A1(_00562_),
    .A2(_03999_),
    .ZN(_04014_));
 OAI21_X1 _20547_ (.A(_04014_),
    .B1(_03669_),
    .B2(_03817_),
    .ZN(_04015_));
 AOI22_X2 _20548_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(_03986_),
    .B1(_04015_),
    .B2(_03990_),
    .ZN(_14192_));
 INV_X1 _20549_ (.A(_15624_),
    .ZN(_14200_));
 NAND2_X1 _20550_ (.A1(_03695_),
    .A2(_03703_),
    .ZN(_14210_));
 OR2_X1 _20551_ (.A1(_00563_),
    .A2(_03999_),
    .ZN(_04016_));
 OAI21_X1 _20552_ (.A(_04016_),
    .B1(_03669_),
    .B2(_03819_),
    .ZN(_04017_));
 AOI22_X2 _20553_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_03658_),
    .B1(_04017_),
    .B2(_11431_),
    .ZN(_14223_));
 NAND2_X1 _20554_ (.A1(_03683_),
    .A2(_03729_),
    .ZN(_14245_));
 NAND2_X1 _20555_ (.A1(_03702_),
    .A2(_03703_),
    .ZN(_14250_));
 NOR2_X1 _20556_ (.A1(_03821_),
    .A2(_03669_),
    .ZN(_04018_));
 AOI21_X1 _20557_ (.A(_04018_),
    .B1(_03988_),
    .B2(_00564_),
    .ZN(_04019_));
 AOI22_X2 _20558_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(_03658_),
    .B1(_04019_),
    .B2(_11431_),
    .ZN(_14263_));
 NAND2_X1 _20559_ (.A1(_03690_),
    .A2(_03729_),
    .ZN(_14285_));
 NAND2_X1 _20560_ (.A1(_03994_),
    .A2(_03708_),
    .ZN(_14290_));
 OR2_X1 _20561_ (.A1(_00565_),
    .A2(_03999_),
    .ZN(_04020_));
 OAI21_X1 _20562_ (.A(_04020_),
    .B1(_03669_),
    .B2(_03824_),
    .ZN(_04021_));
 AOI22_X2 _20563_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(_03658_),
    .B1(_04021_),
    .B2(_11431_),
    .ZN(_14306_));
 NAND2_X1 _20564_ (.A1(_03702_),
    .A2(net336),
    .ZN(_14328_));
 NAND2_X1 _20565_ (.A1(_03994_),
    .A2(_03715_),
    .ZN(_14333_));
 NAND2_X1 _20566_ (.A1(_03702_),
    .A2(_03729_),
    .ZN(_14379_));
 NAND2_X1 _20567_ (.A1(net325),
    .A2(_03735_),
    .ZN(_14387_));
 NOR2_X1 _20568_ (.A1(_03829_),
    .A2(_03669_),
    .ZN(_04022_));
 BUF_X2 _20569_ (.A(_00597_),
    .Z(_04023_));
 AOI21_X1 _20570_ (.A(_04022_),
    .B1(_03988_),
    .B2(_04023_),
    .ZN(_04024_));
 AOI22_X2 _20571_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(_03658_),
    .B1(_04024_),
    .B2(_11431_),
    .ZN(_14408_));
 NAND2_X1 _20572_ (.A1(_03715_),
    .A2(net336),
    .ZN(_14435_));
 NAND2_X1 _20573_ (.A1(net325),
    .A2(_03742_),
    .ZN(_14443_));
 NOR2_X1 _20574_ (.A1(_03831_),
    .A2(_11433_),
    .ZN(_04025_));
 BUF_X2 _20575_ (.A(_00628_),
    .Z(_04026_));
 AOI21_X1 _20576_ (.A(_04025_),
    .B1(_03988_),
    .B2(_04026_),
    .ZN(_04027_));
 AOI22_X2 _20577_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_03658_),
    .B1(_04027_),
    .B2(_11431_),
    .ZN(_14463_));
 NAND2_X4 _20578_ (.A1(_03998_),
    .A2(_03749_),
    .ZN(_14501_));
 NAND2_X1 _20579_ (.A1(_03683_),
    .A2(_03774_),
    .ZN(_14541_));
 NAND2_X1 _20580_ (.A1(_03995_),
    .A2(_03735_),
    .ZN(_14555_));
 NAND2_X1 _20581_ (.A1(net323),
    .A2(_03749_),
    .ZN(_14567_));
 NAND2_X1 _20582_ (.A1(_03695_),
    .A2(_03765_),
    .ZN(_14611_));
 NAND2_X1 _20583_ (.A1(_03697_),
    .A2(_03763_),
    .ZN(_14635_));
 NAND2_X1 _20584_ (.A1(_03995_),
    .A2(net431),
    .ZN(_14684_));
 NAND2_X1 _20585_ (.A1(net337),
    .A2(_03755_),
    .ZN(_14742_));
 NAND2_X1 _20586_ (.A1(_03715_),
    .A2(_03765_),
    .ZN(_14787_));
 NAND2_X1 _20587_ (.A1(_03697_),
    .A2(_03812_),
    .ZN(_14810_));
 NAND2_X1 _20588_ (.A1(_03715_),
    .A2(_03774_),
    .ZN(_14844_));
 NAND2_X1 _20589_ (.A1(net337),
    .A2(_03770_),
    .ZN(_14857_));
 NAND2_X1 _20590_ (.A1(net324),
    .A2(_03812_),
    .ZN(_14867_));
 NAND2_X1 _20591_ (.A1(net337),
    .A2(_03776_),
    .ZN(_14910_));
 NAND2_X1 _20592_ (.A1(_03742_),
    .A2(_03765_),
    .ZN(_14951_));
 NAND2_X1 _20593_ (.A1(_03826_),
    .A2(_03755_),
    .ZN(_14956_));
 NAND2_X1 _20594_ (.A1(_03742_),
    .A2(_03774_),
    .ZN(_15004_));
 INV_X1 _20595_ (.A(_14816_),
    .ZN(_14817_));
 NAND2_X1 _20596_ (.A1(_03826_),
    .A2(_03770_),
    .ZN(_15055_));
 NAND2_X1 _20597_ (.A1(net291),
    .A2(_03770_),
    .ZN(_15137_));
 NAND2_X1 _20598_ (.A1(net291),
    .A2(_03776_),
    .ZN(_15176_));
 NAND2_X1 _20599_ (.A1(net291),
    .A2(_03784_),
    .ZN(_15213_));
 NAND2_X1 _20600_ (.A1(_03996_),
    .A2(_03784_),
    .ZN(_15252_));
 INV_X2 _20601_ (.A(_15023_),
    .ZN(_15068_));
 NAND2_X1 _20602_ (.A1(_03996_),
    .A2(_03798_),
    .ZN(_15291_));
 OR2_X2 _20603_ (.A1(_00137_),
    .A2(_03974_),
    .ZN(_15354_));
 INV_X1 _20604_ (.A(_14186_),
    .ZN(_14187_));
 INV_X1 _20605_ (.A(_14217_),
    .ZN(_14218_));
 INV_X1 _20606_ (.A(_14257_),
    .ZN(_14258_));
 INV_X1 _20607_ (.A(_14278_),
    .ZN(_14280_));
 INV_X1 _20608_ (.A(_14297_),
    .ZN(_14298_));
 INV_X2 _20609_ (.A(_14321_),
    .ZN(_14323_));
 INV_X1 _20610_ (.A(_14340_),
    .ZN(_14341_));
 INV_X1 _20611_ (.A(_14367_),
    .ZN(_14368_));
 INV_X1 _20612_ (.A(_14394_),
    .ZN(_14395_));
 INV_X1 _20613_ (.A(_14405_),
    .ZN(_14419_));
 INV_X1 _20614_ (.A(_14418_),
    .ZN(_14420_));
 INV_X2 _20615_ (.A(_14450_),
    .ZN(_14451_));
 INV_X2 _20616_ (.A(_14460_),
    .ZN(_14474_));
 INV_X1 _20617_ (.A(_14473_),
    .ZN(_14475_));
 INV_X1 _20618_ (.A(_14508_),
    .ZN(_14509_));
 INV_X2 _20619_ (.A(_14517_),
    .ZN(_14531_));
 INV_X1 _20620_ (.A(_14530_),
    .ZN(_14532_));
 INV_X1 _20621_ (.A(_14564_),
    .ZN(_14580_));
 INV_X1 _20622_ (.A(_14574_),
    .ZN(_14575_));
 INV_X1 _20623_ (.A(_14588_),
    .ZN(_14590_));
 INV_X1 _20624_ (.A(_14601_),
    .ZN(_14603_));
 INV_X1 _20625_ (.A(_14618_),
    .ZN(_14619_));
 INV_X1 _20626_ (.A(_14642_),
    .ZN(_14643_));
 INV_X1 _20627_ (.A(_14654_),
    .ZN(_14656_));
 INV_X1 _20628_ (.A(_14678_),
    .ZN(_14679_));
 INV_X1 _20629_ (.A(_14701_),
    .ZN(_14702_));
 INV_X1 _20630_ (.A(_14711_),
    .ZN(_14712_));
 INV_X1 _20631_ (.A(_14721_),
    .ZN(_14722_));
 INV_X1 _20632_ (.A(_14736_),
    .ZN(_14737_));
 INV_X1 _20633_ (.A(_14768_),
    .ZN(_14769_));
 INV_X1 _20634_ (.A(_14778_),
    .ZN(_14779_));
 INV_X1 _20635_ (.A(_14794_),
    .ZN(_14795_));
 INV_X1 _20636_ (.A(_14826_),
    .ZN(_14827_));
 INV_X1 _20637_ (.A(_14835_),
    .ZN(_14836_));
 INV_X1 _20638_ (.A(_14851_),
    .ZN(_14852_));
 INV_X1 _20639_ (.A(_14878_),
    .ZN(_14879_));
 INV_X1 _20640_ (.A(_14888_),
    .ZN(_14889_));
 INV_X1 _20641_ (.A(_14904_),
    .ZN(_14905_));
 INV_X1 _20642_ (.A(_14925_),
    .ZN(_14926_));
 INV_X1 _20643_ (.A(_14933_),
    .ZN(_14934_));
 INV_X1 _20644_ (.A(_14942_),
    .ZN(_14943_));
 INV_X1 _20645_ (.A(_14986_),
    .ZN(_14988_));
 INV_X1 _20646_ (.A(_14995_),
    .ZN(_14996_));
 INV_X1 _20647_ (.A(_15032_),
    .ZN(_15034_));
 INV_X1 _20648_ (.A(_15041_),
    .ZN(_15042_));
 INV_X1 _20649_ (.A(_15075_),
    .ZN(_15077_));
 INV_X1 _20650_ (.A(_15084_),
    .ZN(_15085_));
 INV_X2 _20651_ (.A(_15107_),
    .ZN(_15108_));
 INV_X1 _20652_ (.A(_15119_),
    .ZN(_15120_));
 INV_X1 _20653_ (.A(_15128_),
    .ZN(_15129_));
 INV_X1 _20654_ (.A(_15158_),
    .ZN(_15159_));
 INV_X1 _20655_ (.A(_15167_),
    .ZN(_15168_));
 INV_X1 _20656_ (.A(_15195_),
    .ZN(_15196_));
 INV_X1 _20657_ (.A(_15204_),
    .ZN(_15205_));
 INV_X1 _20658_ (.A(_15234_),
    .ZN(_15235_));
 INV_X1 _20659_ (.A(_15243_),
    .ZN(_15244_));
 INV_X1 _20660_ (.A(_15258_),
    .ZN(_15262_));
 INV_X1 _20661_ (.A(_15268_),
    .ZN(_15269_));
 INV_X1 _20662_ (.A(_15274_),
    .ZN(_15275_));
 INV_X1 _20663_ (.A(_15283_),
    .ZN(_15284_));
 INV_X1 _20664_ (.A(_15297_),
    .ZN(_15298_));
 INV_X1 _20665_ (.A(_15304_),
    .ZN(_15305_));
 INV_X1 _20666_ (.A(_15310_),
    .ZN(_15311_));
 INV_X1 _20667_ (.A(_15318_),
    .ZN(_15319_));
 INV_X1 _20668_ (.A(_15333_),
    .ZN(_15334_));
 INV_X1 _20669_ (.A(_15341_),
    .ZN(_15824_));
 INV_X1 _20670_ (.A(_15345_),
    .ZN(_15346_));
 INV_X1 _20671_ (.A(_14087_),
    .ZN(_14114_));
 INV_X1 _20672_ (.A(_14107_),
    .ZN(_14137_));
 INV_X1 _20673_ (.A(_14130_),
    .ZN(_14164_));
 INV_X1 _20674_ (.A(_14153_),
    .ZN(_14195_));
 INV_X1 _20675_ (.A(_14185_),
    .ZN(_14226_));
 INV_X1 _20676_ (.A(_14216_),
    .ZN(_14266_));
 INV_X1 _20677_ (.A(_14237_),
    .ZN(_14279_));
 INV_X1 _20678_ (.A(_14256_),
    .ZN(_14309_));
 INV_X1 _20679_ (.A(_14277_),
    .ZN(_14322_));
 INV_X1 _20680_ (.A(_14296_),
    .ZN(_14357_));
 INV_X1 _20681_ (.A(_14320_),
    .ZN(_14369_));
 INV_X1 _20682_ (.A(_14339_),
    .ZN(_14411_));
 INV_X1 _20683_ (.A(_14350_),
    .ZN(_14421_));
 INV_X1 _20684_ (.A(_14363_),
    .ZN(_14425_));
 INV_X1 _20685_ (.A(_14366_),
    .ZN(_14424_));
 INV_X1 _20686_ (.A(_14375_),
    .ZN(_14438_));
 INV_X1 _20687_ (.A(_14393_),
    .ZN(_14466_));
 INV_X1 _20688_ (.A(_14404_),
    .ZN(_14476_));
 INV_X1 _20689_ (.A(_14417_),
    .ZN(_14479_));
 INV_X1 _20690_ (.A(_14449_),
    .ZN(_14523_));
 INV_X1 _20691_ (.A(_14459_),
    .ZN(_14533_));
 INV_X1 _20692_ (.A(_14472_),
    .ZN(_14536_));
 INV_X1 _20693_ (.A(_14485_),
    .ZN(_14558_));
 INV_X1 _20694_ (.A(_14497_),
    .ZN(_14581_));
 INV_X1 _20695_ (.A(_14507_),
    .ZN(_14589_));
 INV_X1 _20696_ (.A(_14516_),
    .ZN(_14602_));
 INV_X1 _20697_ (.A(_14529_),
    .ZN(_14606_));
 INV_X1 _20698_ (.A(_14547_),
    .ZN(_14627_));
 INV_X1 _20699_ (.A(_14551_),
    .ZN(_14630_));
 INV_X1 _20700_ (.A(_14563_),
    .ZN(_14648_));
 INV_X1 _20701_ (.A(_14573_),
    .ZN(_14655_));
 INV_X1 _20702_ (.A(_14587_),
    .ZN(_14657_));
 INV_X1 _20703_ (.A(_14596_),
    .ZN(_14661_));
 INV_X1 _20704_ (.A(_14600_),
    .ZN(_14666_));
 INV_X1 _20705_ (.A(_14617_),
    .ZN(_14687_));
 INV_X1 _20706_ (.A(_14641_),
    .ZN(_14714_));
 INV_X1 _20707_ (.A(_14653_),
    .ZN(_14713_));
 INV_X1 _20708_ (.A(_14677_),
    .ZN(_14745_));
 INV_X1 _20709_ (.A(_14700_),
    .ZN(_14770_));
 INV_X1 _20710_ (.A(_14710_),
    .ZN(_14771_));
 INV_X1 _20711_ (.A(_14720_),
    .ZN(_14782_));
 INV_X1 _20712_ (.A(_14735_),
    .ZN(_14803_));
 INV_X1 _20713_ (.A(_14767_),
    .ZN(_14828_));
 INV_X1 _20714_ (.A(_14777_),
    .ZN(_14839_));
 INV_X1 _20715_ (.A(_14793_),
    .ZN(_14860_));
 INV_X1 _20716_ (.A(_14825_),
    .ZN(_14881_));
 INV_X1 _20717_ (.A(_14834_),
    .ZN(_14892_));
 INV_X1 _20718_ (.A(_14850_),
    .ZN(_14913_));
 INV_X1 _20719_ (.A(_14877_),
    .ZN(_14935_));
 INV_X1 _20720_ (.A(_14887_),
    .ZN(_14946_));
 INV_X1 _20721_ (.A(_14903_),
    .ZN(_14966_));
 INV_X1 _20722_ (.A(_14924_),
    .ZN(_14979_));
 INV_X1 _20723_ (.A(_14932_),
    .ZN(_14987_));
 INV_X1 _20724_ (.A(_14941_),
    .ZN(_14999_));
 INV_X1 _20725_ (.A(_14985_),
    .ZN(_15033_));
 INV_X1 _20726_ (.A(_14994_),
    .ZN(_15045_));
 INV_X1 _20727_ (.A(_15031_),
    .ZN(_15076_));
 INV_X1 _20728_ (.A(_15040_),
    .ZN(_15088_));
 INV_X1 _20729_ (.A(_15074_),
    .ZN(_15121_));
 INV_X1 _20730_ (.A(_15083_),
    .ZN(_15132_));
 INV_X2 _20731_ (.A(_15106_),
    .ZN(_15147_));
 INV_X1 _20732_ (.A(_15118_),
    .ZN(_15160_));
 INV_X1 _20733_ (.A(_15127_),
    .ZN(_15171_));
 INV_X1 _20734_ (.A(_15157_),
    .ZN(_15197_));
 INV_X1 _20735_ (.A(_15166_),
    .ZN(_15208_));
 INV_X1 _20736_ (.A(_15194_),
    .ZN(_15236_));
 INV_X1 _20737_ (.A(_15203_),
    .ZN(_15247_));
 INV_X1 _20738_ (.A(_15219_),
    .ZN(_15259_));
 INV_X1 _20739_ (.A(_15233_),
    .ZN(_15276_));
 INV_X1 _20740_ (.A(_15242_),
    .ZN(_15287_));
 INV_X1 _20741_ (.A(_15257_),
    .ZN(_15299_));
 INV_X1 _20742_ (.A(_15273_),
    .ZN(_15312_));
 INV_X1 _20743_ (.A(_15282_),
    .ZN(_15322_));
 INV_X1 _20744_ (.A(_15317_),
    .ZN(_15349_));
 CLKBUF_X3 _20745_ (.A(_03449_),
    .Z(_04028_));
 CLKBUF_X3 _20746_ (.A(_04028_),
    .Z(_04029_));
 BUF_X8 _20747_ (.A(_12099_),
    .Z(_04030_));
 XNOR2_X1 _20748_ (.A(_15834_),
    .B(_04030_),
    .ZN(_04031_));
 NOR2_X1 _20749_ (.A1(_04029_),
    .A2(_04031_),
    .ZN(_04032_));
 BUF_X4 _20750_ (.A(_03405_),
    .Z(_04033_));
 CLKBUF_X3 _20751_ (.A(_04033_),
    .Z(_04034_));
 CLKBUF_X3 _20752_ (.A(_03406_),
    .Z(_04035_));
 OAI22_X1 _20753_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_03675_),
    .ZN(_04036_));
 BUF_X4 _20754_ (.A(_03407_),
    .Z(_04037_));
 BUF_X4 _20755_ (.A(_03402_),
    .Z(_04038_));
 OAI22_X1 _20756_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_04037_),
    .B1(_03681_),
    .B2(_04038_),
    .ZN(_04039_));
 CLKBUF_X3 _20757_ (.A(_03406_),
    .Z(_04040_));
 CLKBUF_X3 _20758_ (.A(_04040_),
    .Z(_04041_));
 AOI21_X1 _20759_ (.A(_04036_),
    .B1(_04039_),
    .B2(_04041_),
    .ZN(_04042_));
 BUF_X4 _20760_ (.A(_04028_),
    .Z(_04043_));
 AOI21_X2 _20761_ (.A(_04032_),
    .B1(_04042_),
    .B2(_04043_),
    .ZN(_15369_));
 BUF_X4 _20762_ (.A(_03407_),
    .Z(_04044_));
 OR2_X2 _20763_ (.A1(_10777_),
    .A2(_10812_),
    .ZN(_04045_));
 OAI221_X1 _20764_ (.A(_03406_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B2(_04044_),
    .C1(_04038_),
    .C2(_04045_),
    .ZN(_04046_));
 OAI21_X1 _20765_ (.A(_04046_),
    .B1(_04040_),
    .B2(_03660_),
    .ZN(_04047_));
 BUF_X2 _20766_ (.A(_04034_),
    .Z(_04048_));
 OAI21_X1 _20767_ (.A(_04047_),
    .B1(_04048_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .ZN(_04049_));
 BUF_X16 _20768_ (.A(_04030_),
    .Z(_04050_));
 XNOR2_X2 _20769_ (.A(_15835_),
    .B(_04050_),
    .ZN(_04051_));
 BUF_X2 _20770_ (.A(_11409_),
    .Z(_04052_));
 MUX2_X1 _20771_ (.A(_04049_),
    .B(_04051_),
    .S(_04052_),
    .Z(_14065_));
 XNOR2_X1 _20772_ (.A(_15857_),
    .B(_04050_),
    .ZN(_04053_));
 BUF_X4 _20773_ (.A(_04033_),
    .Z(_04054_));
 BUF_X4 _20774_ (.A(_03402_),
    .Z(_04055_));
 OAI222_X2 _20775_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .B2(_04054_),
    .C1(net294),
    .C2(_04055_),
    .ZN(_04056_));
 MUX2_X1 _20776_ (.A(_10972_),
    .B(_04056_),
    .S(_04040_),
    .Z(_04057_));
 CLKBUF_X3 _20777_ (.A(_04028_),
    .Z(_04058_));
 MUX2_X1 _20778_ (.A(_04053_),
    .B(_04057_),
    .S(_04058_),
    .Z(_15375_));
 XNOR2_X1 _20779_ (.A(_15860_),
    .B(_04030_),
    .ZN(_04059_));
 NOR2_X1 _20780_ (.A1(_04029_),
    .A2(_04059_),
    .ZN(_04060_));
 OAI22_X1 _20781_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_11019_),
    .ZN(_04061_));
 OAI22_X1 _20782_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .B1(net319),
    .B2(_04038_),
    .ZN(_04062_));
 AOI21_X1 _20783_ (.A(_04061_),
    .B1(_04062_),
    .B2(_04041_),
    .ZN(_04063_));
 AOI21_X1 _20784_ (.A(_04060_),
    .B1(_04063_),
    .B2(_04043_),
    .ZN(_15379_));
 XNOR2_X1 _20785_ (.A(_15873_),
    .B(_04050_),
    .ZN(_04064_));
 OAI222_X2 _20786_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .B2(_04054_),
    .C1(_11591_),
    .C2(_04055_),
    .ZN(_04065_));
 MUX2_X1 _20787_ (.A(_11057_),
    .B(_04065_),
    .S(_04040_),
    .Z(_04066_));
 MUX2_X1 _20788_ (.A(_04064_),
    .B(_04066_),
    .S(_04058_),
    .Z(_15383_));
 XNOR2_X1 _20789_ (.A(_15880_),
    .B(net296),
    .ZN(_04067_));
 OAI222_X2 _20790_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .B2(_04033_),
    .C1(_11629_),
    .C2(_04055_),
    .ZN(_04068_));
 MUX2_X1 _20791_ (.A(_11115_),
    .B(_04068_),
    .S(_04040_),
    .Z(_04069_));
 MUX2_X1 _20792_ (.A(_04067_),
    .B(_04069_),
    .S(_04058_),
    .Z(_15387_));
 XNOR2_X1 _20793_ (.A(_15888_),
    .B(net296),
    .ZN(_04070_));
 AND3_X1 _20794_ (.A1(_03401_),
    .A2(_03402_),
    .A3(_04033_),
    .ZN(_04071_));
 OAI222_X2 _20795_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .B2(_04033_),
    .C1(_11672_),
    .C2(_03402_),
    .ZN(_04072_));
 NOR2_X1 _20796_ (.A1(_04071_),
    .A2(_04072_),
    .ZN(_04073_));
 AOI21_X1 _20797_ (.A(_04073_),
    .B1(_04071_),
    .B2(_11158_),
    .ZN(_04074_));
 MUX2_X1 _20798_ (.A(_04070_),
    .B(_04074_),
    .S(_04058_),
    .Z(_15391_));
 OR3_X1 _20799_ (.A1(_00561_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04075_));
 OAI21_X1 _20800_ (.A(_04075_),
    .B1(_15897_),
    .B2(_04043_),
    .ZN(_15395_));
 OAI221_X1 _20801_ (.A(_03406_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B2(_03407_),
    .C1(_04038_),
    .C2(_03732_),
    .ZN(_04076_));
 OAI21_X1 _20802_ (.A(_04076_),
    .B1(_04040_),
    .B2(_11241_),
    .ZN(_04077_));
 OAI21_X1 _20803_ (.A(_04077_),
    .B1(_04048_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .ZN(_04078_));
 XNOR2_X1 _20804_ (.A(_15904_),
    .B(net317),
    .ZN(_04079_));
 MUX2_X1 _20805_ (.A(_04078_),
    .B(_04079_),
    .S(_04052_),
    .Z(_15399_));
 XNOR2_X1 _20806_ (.A(_15908_),
    .B(_11863_),
    .ZN(_04080_));
 OAI222_X2 _20807_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .B2(_04033_),
    .C1(_11824_),
    .C2(_04055_),
    .ZN(_04081_));
 MUX2_X1 _20808_ (.A(_11279_),
    .B(_04081_),
    .S(_03406_),
    .Z(_04082_));
 MUX2_X1 _20809_ (.A(_04080_),
    .B(_04082_),
    .S(_04058_),
    .Z(_15403_));
 OAI221_X1 _20810_ (.A(_03406_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B2(_03407_),
    .C1(_04038_),
    .C2(_11898_),
    .ZN(_04083_));
 OAI21_X1 _20811_ (.A(_04083_),
    .B1(_04040_),
    .B2(_11313_),
    .ZN(_04084_));
 OAI21_X1 _20812_ (.A(_04084_),
    .B1(_04048_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .ZN(_04085_));
 XNOR2_X1 _20813_ (.A(_15920_),
    .B(net317),
    .ZN(_04086_));
 MUX2_X1 _20814_ (.A(_04085_),
    .B(_04086_),
    .S(_04052_),
    .Z(_15407_));
 OR3_X1 _20815_ (.A1(_00565_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04087_));
 OAI21_X1 _20816_ (.A(_04087_),
    .B1(_04043_),
    .B2(_15928_),
    .ZN(_15411_));
 OR3_X1 _20817_ (.A1(_00566_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04088_));
 OAI21_X1 _20818_ (.A(_04088_),
    .B1(_04043_),
    .B2(_15936_),
    .ZN(_15415_));
 OR3_X1 _20819_ (.A1(_04023_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04089_));
 CLKBUF_X3 _20820_ (.A(_04028_),
    .Z(_04090_));
 OAI21_X1 _20821_ (.A(_04089_),
    .B1(_15944_),
    .B2(_04090_),
    .ZN(_15419_));
 XNOR2_X1 _20822_ (.A(net296),
    .B(_15953_),
    .ZN(_04091_));
 NOR2_X1 _20823_ (.A1(_04029_),
    .A2(_04091_),
    .ZN(_04092_));
 OAI22_X2 _20824_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_12144_),
    .ZN(_04093_));
 OAI22_X2 _20825_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B1(_12177_),
    .B2(_04038_),
    .ZN(_04094_));
 AOI21_X2 _20826_ (.A(_04093_),
    .B1(_04094_),
    .B2(_04041_),
    .ZN(_04095_));
 AOI21_X2 _20827_ (.A(_04092_),
    .B1(_04095_),
    .B2(_04043_),
    .ZN(_15423_));
 XNOR2_X1 _20828_ (.A(net296),
    .B(_15956_),
    .ZN(_04096_));
 NOR2_X1 _20829_ (.A1(_04029_),
    .A2(_04096_),
    .ZN(_04097_));
 OAI22_X1 _20830_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_12221_),
    .ZN(_04098_));
 OAI22_X1 _20831_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .B1(_12254_),
    .B2(_04038_),
    .ZN(_04099_));
 AOI21_X1 _20832_ (.A(_04098_),
    .B1(_04099_),
    .B2(_04041_),
    .ZN(_04100_));
 AOI21_X2 _20833_ (.A(_04097_),
    .B1(_04100_),
    .B2(_04043_),
    .ZN(_15427_));
 XNOR2_X1 _20834_ (.A(net296),
    .B(_15969_),
    .ZN(_04101_));
 NOR2_X1 _20835_ (.A1(_04058_),
    .A2(_04101_),
    .ZN(_04102_));
 OAI22_X1 _20836_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_12316_),
    .ZN(_04103_));
 OAI22_X1 _20837_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B1(_12350_),
    .B2(_04038_),
    .ZN(_04104_));
 AOI21_X1 _20838_ (.A(_04103_),
    .B1(_04104_),
    .B2(_04041_),
    .ZN(_04105_));
 AOI21_X2 _20839_ (.A(_04102_),
    .B1(_04105_),
    .B2(_04043_),
    .ZN(_15431_));
 XNOR2_X1 _20840_ (.A(net317),
    .B(_15977_),
    .ZN(_04106_));
 BUF_X4 _20841_ (.A(_04033_),
    .Z(_04107_));
 OAI222_X2 _20842_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .B2(_04107_),
    .C1(_12425_),
    .C2(_04038_),
    .ZN(_04108_));
 NAND2_X1 _20843_ (.A1(_04035_),
    .A2(_04108_),
    .ZN(_04109_));
 OAI21_X1 _20844_ (.A(_04109_),
    .B1(_04041_),
    .B2(_12392_),
    .ZN(_04110_));
 MUX2_X1 _20845_ (.A(_04106_),
    .B(_04110_),
    .S(_04058_),
    .Z(_15435_));
 XNOR2_X1 _20846_ (.A(net317),
    .B(_15980_),
    .ZN(_04111_));
 BUF_X4 _20847_ (.A(_03402_),
    .Z(_04112_));
 OAI222_X2 _20848_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .B2(_04107_),
    .C1(_12514_),
    .C2(_04112_),
    .ZN(_04113_));
 NAND2_X1 _20849_ (.A1(_04035_),
    .A2(_04113_),
    .ZN(_04114_));
 OAI21_X1 _20850_ (.A(_04114_),
    .B1(_04041_),
    .B2(net347),
    .ZN(_04115_));
 MUX2_X1 _20851_ (.A(_04111_),
    .B(_04115_),
    .S(_04058_),
    .Z(_15439_));
 OR3_X1 _20852_ (.A1(_00783_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04116_));
 OAI21_X1 _20853_ (.A(_04116_),
    .B1(_15992_),
    .B2(_04090_),
    .ZN(_15443_));
 CLKBUF_X3 _20854_ (.A(_11863_),
    .Z(_04117_));
 XNOR2_X1 _20855_ (.A(_04117_),
    .B(_16000_),
    .ZN(_04118_));
 OAI222_X2 _20856_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .B2(_04107_),
    .C1(net358),
    .C2(_04112_),
    .ZN(_04119_));
 NAND2_X1 _20857_ (.A1(_04035_),
    .A2(_04119_),
    .ZN(_04120_));
 OAI21_X1 _20858_ (.A(_04120_),
    .B1(_04041_),
    .B2(_12651_),
    .ZN(_04121_));
 MUX2_X1 _20859_ (.A(_04118_),
    .B(_04121_),
    .S(_04058_),
    .Z(_15447_));
 OR3_X1 _20860_ (.A1(_00845_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04122_));
 OAI21_X1 _20861_ (.A(_04122_),
    .B1(_16005_),
    .B2(_04090_),
    .ZN(_15451_));
 XNOR2_X1 _20862_ (.A(_04117_),
    .B(_16016_),
    .ZN(_04123_));
 OAI222_X2 _20863_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .B2(_04107_),
    .C1(_03713_),
    .C2(_04112_),
    .ZN(_04124_));
 NAND2_X1 _20864_ (.A1(_04035_),
    .A2(_04124_),
    .ZN(_04125_));
 OAI21_X1 _20865_ (.A(_04125_),
    .B1(_04041_),
    .B2(_12823_),
    .ZN(_04126_));
 MUX2_X1 _20866_ (.A(_04123_),
    .B(_04126_),
    .S(_04058_),
    .Z(_15455_));
 XNOR2_X1 _20867_ (.A(_04117_),
    .B(_16021_),
    .ZN(_04127_));
 BUF_X2 _20868_ (.A(_03406_),
    .Z(_04128_));
 OAI222_X2 _20869_ (.A1(_04037_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .B2(_04107_),
    .C1(_03724_),
    .C2(_04112_),
    .ZN(_04129_));
 NAND2_X1 _20870_ (.A1(_04128_),
    .A2(_04129_),
    .ZN(_04130_));
 OAI21_X1 _20871_ (.A(_04130_),
    .B1(_04041_),
    .B2(net421),
    .ZN(_04131_));
 CLKBUF_X3 _20872_ (.A(_04028_),
    .Z(_04132_));
 MUX2_X1 _20873_ (.A(_04127_),
    .B(_04131_),
    .S(_04132_),
    .Z(_15459_));
 OR3_X1 _20874_ (.A1(_03817_),
    .A2(_04052_),
    .A3(_04048_),
    .ZN(_04133_));
 OAI21_X1 _20875_ (.A(_04133_),
    .B1(_16029_),
    .B2(_04090_),
    .ZN(_15463_));
 CLKBUF_X2 _20876_ (.A(_11409_),
    .Z(_04134_));
 CLKBUF_X2 _20877_ (.A(_04107_),
    .Z(_04135_));
 OR3_X1 _20878_ (.A1(_03819_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04136_));
 OAI21_X1 _20879_ (.A(_04136_),
    .B1(_16040_),
    .B2(_04090_),
    .ZN(_15467_));
 XNOR2_X1 _20880_ (.A(_04117_),
    .B(_16048_),
    .ZN(_04137_));
 BUF_X4 _20881_ (.A(_03407_),
    .Z(_04138_));
 OAI222_X2 _20882_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .B2(_04107_),
    .C1(net352),
    .C2(_04112_),
    .ZN(_04139_));
 NAND2_X1 _20883_ (.A1(_04128_),
    .A2(_04139_),
    .ZN(_04140_));
 BUF_X2 _20884_ (.A(_04040_),
    .Z(_04141_));
 OAI21_X1 _20885_ (.A(_04140_),
    .B1(_04141_),
    .B2(_13155_),
    .ZN(_04142_));
 MUX2_X1 _20886_ (.A(_04137_),
    .B(_04142_),
    .S(_04132_),
    .Z(_15471_));
 XNOR2_X1 _20887_ (.A(_04117_),
    .B(_16053_),
    .ZN(_04143_));
 OAI222_X2 _20888_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .B2(_04107_),
    .C1(net342),
    .C2(_04112_),
    .ZN(_04144_));
 NAND2_X1 _20889_ (.A1(_04128_),
    .A2(_04144_),
    .ZN(_04145_));
 OAI21_X1 _20890_ (.A(_04145_),
    .B1(_04141_),
    .B2(_13224_),
    .ZN(_04146_));
 MUX2_X1 _20891_ (.A(_04143_),
    .B(_04146_),
    .S(_04132_),
    .Z(_15475_));
 OR3_X1 _20892_ (.A1(_03827_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04147_));
 OAI21_X1 _20893_ (.A(_04147_),
    .B1(_16064_),
    .B2(_04090_),
    .ZN(_15479_));
 XNOR2_X1 _20894_ (.A(_04117_),
    .B(_16069_),
    .ZN(_04148_));
 OAI222_X2 _20895_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .B2(_04107_),
    .C1(_03769_),
    .C2(_04112_),
    .ZN(_04149_));
 NAND2_X1 _20896_ (.A1(_04128_),
    .A2(_04149_),
    .ZN(_04150_));
 OAI21_X1 _20897_ (.A(_04150_),
    .B1(_04141_),
    .B2(_03166_),
    .ZN(_04151_));
 MUX2_X1 _20898_ (.A(_04148_),
    .B(_04151_),
    .S(_04132_),
    .Z(_15483_));
 OR3_X1 _20899_ (.A1(_01124_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04152_));
 OAI21_X1 _20900_ (.A(_04152_),
    .B1(_16080_),
    .B2(_04090_),
    .ZN(_15487_));
 INV_X1 _20901_ (.A(_15495_),
    .ZN(_15491_));
 NOR2_X1 _20902_ (.A1(_10920_),
    .A2(_15912_),
    .ZN(_15499_));
 INV_X1 _20903_ (.A(_15904_),
    .ZN(_15900_));
 NAND2_X1 _20904_ (.A1(_10922_),
    .A2(_15900_),
    .ZN(_15503_));
 INV_X1 _20905_ (.A(_14078_),
    .ZN(_15557_));
 INV_X1 _20906_ (.A(_14116_),
    .ZN(_15592_));
 INV_X1 _20907_ (.A(_14121_),
    .ZN(_14122_));
 INV_X1 _20908_ (.A(_14139_),
    .ZN(_15608_));
 INV_X1 _20909_ (.A(_14115_),
    .ZN(_15609_));
 INV_X1 _20910_ (.A(_14144_),
    .ZN(_15616_));
 INV_X1 _20911_ (.A(_14166_),
    .ZN(_15622_));
 INV_X1 _20912_ (.A(_14171_),
    .ZN(_15626_));
 INV_X1 _20913_ (.A(_14176_),
    .ZN(_15628_));
 INV_X1 _20914_ (.A(_14189_),
    .ZN(_15632_));
 INV_X1 _20915_ (.A(_14197_),
    .ZN(_15637_));
 INV_X1 _20916_ (.A(_14202_),
    .ZN(_15641_));
 INV_X1 _20917_ (.A(_14220_),
    .ZN(_15649_));
 INV_X1 _20918_ (.A(_14228_),
    .ZN(_15653_));
 INV_X1 _20919_ (.A(_14196_),
    .ZN(_15654_));
 INV_X1 _20920_ (.A(_14233_),
    .ZN(_14235_));
 INV_X1 _20921_ (.A(_14247_),
    .ZN(_15659_));
 INV_X1 _20922_ (.A(_14260_),
    .ZN(_15662_));
 INV_X2 _20923_ (.A(_14268_),
    .ZN(_15666_));
 INV_X1 _20924_ (.A(_14227_),
    .ZN(_15667_));
 INV_X1 _20925_ (.A(_14273_),
    .ZN(_14275_));
 INV_X1 _20926_ (.A(_14287_),
    .ZN(_15673_));
 INV_X1 _20927_ (.A(_14303_),
    .ZN(_15679_));
 INV_X2 _20928_ (.A(_14311_),
    .ZN(_15680_));
 INV_X1 _20929_ (.A(_14267_),
    .ZN(_15681_));
 INV_X2 _20930_ (.A(_14316_),
    .ZN(_14318_));
 INV_X1 _20931_ (.A(_14281_),
    .ZN(_15683_));
 INV_X1 _20932_ (.A(_14330_),
    .ZN(_15691_));
 INV_X1 _20933_ (.A(_14346_),
    .ZN(_14349_));
 INV_X1 _20934_ (.A(_14359_),
    .ZN(_15695_));
 INV_X2 _20935_ (.A(_14371_),
    .ZN(_15697_));
 INV_X1 _20936_ (.A(_14400_),
    .ZN(_14403_));
 INV_X1 _20937_ (.A(_14413_),
    .ZN(_15702_));
 INV_X1 _20938_ (.A(_14427_),
    .ZN(_15704_));
 INV_X1 _20939_ (.A(_14440_),
    .ZN(_15711_));
 INV_X1 _20940_ (.A(_14468_),
    .ZN(_15712_));
 INV_X2 _20941_ (.A(_14481_),
    .ZN(_15714_));
 INV_X1 _20942_ (.A(_14493_),
    .ZN(_14496_));
 INV_X1 _20943_ (.A(_14525_),
    .ZN(_15721_));
 INV_X2 _20944_ (.A(_14538_),
    .ZN(_15723_));
 INV_X1 _20945_ (.A(_14543_),
    .ZN(_14549_));
 INV_X1 _20946_ (.A(_14560_),
    .ZN(_14561_));
 INV_X2 _20947_ (.A(_14592_),
    .ZN(_14594_));
 INV_X1 _20948_ (.A(_14512_),
    .ZN(_14598_));
 INV_X1 _20949_ (.A(_14608_),
    .ZN(_15727_));
 INV_X1 _20950_ (.A(_14659_),
    .ZN(_15733_));
 INV_X1 _20951_ (.A(_14668_),
    .ZN(_15736_));
 INV_X1 _20952_ (.A(_14716_),
    .ZN(_15740_));
 INV_X1 _20953_ (.A(_14646_),
    .ZN(_14717_));
 INV_X1 _20954_ (.A(_14726_),
    .ZN(_15742_));
 INV_X1 _20955_ (.A(_14773_),
    .ZN(_15746_));
 INV_X1 _20956_ (.A(_14784_),
    .ZN(_15748_));
 INV_X1 _20957_ (.A(_14830_),
    .ZN(_15752_));
 INV_X1 _20958_ (.A(_14772_),
    .ZN(_15753_));
 INV_X1 _20959_ (.A(_14762_),
    .ZN(_14831_));
 INV_X1 _20960_ (.A(_14783_),
    .ZN(_15754_));
 INV_X1 _20961_ (.A(_14883_),
    .ZN(_15758_));
 INV_X1 _20962_ (.A(_14894_),
    .ZN(_15760_));
 INV_X1 _20963_ (.A(_14868_),
    .ZN(_14922_));
 INV_X1 _20964_ (.A(_14937_),
    .ZN(_15764_));
 INV_X1 _20965_ (.A(_14882_),
    .ZN(_15765_));
 INV_X1 _20966_ (.A(_14872_),
    .ZN(_14938_));
 INV_X1 _20967_ (.A(_14893_),
    .ZN(_15766_));
 INV_X1 _20968_ (.A(_14990_),
    .ZN(_15770_));
 INV_X1 _20969_ (.A(_14927_),
    .ZN(_14991_));
 INV_X1 _20970_ (.A(_15001_),
    .ZN(_15772_));
 INV_X1 _20971_ (.A(_15036_),
    .ZN(_15776_));
 INV_X1 _20972_ (.A(_14989_),
    .ZN(_15777_));
 INV_X1 _20973_ (.A(_15000_),
    .ZN(_15778_));
 INV_X1 _20974_ (.A(_15035_),
    .ZN(_15782_));
 INV_X1 _20975_ (.A(_15026_),
    .ZN(_15081_));
 INV_X1 _20976_ (.A(_15090_),
    .ZN(_15784_));
 INV_X1 _20977_ (.A(_15123_),
    .ZN(_15788_));
 INV_X1 _20978_ (.A(_15069_),
    .ZN(_15125_));
 INV_X1 _20979_ (.A(_15134_),
    .ZN(_15790_));
 INV_X1 _20980_ (.A(_15162_),
    .ZN(_15794_));
 INV_X1 _20981_ (.A(_15122_),
    .ZN(_15795_));
 INV_X1 _20982_ (.A(_15113_),
    .ZN(_15163_));
 INV_X1 _20983_ (.A(_15133_),
    .ZN(_15796_));
 INV_X1 _20984_ (.A(_15199_),
    .ZN(_15800_));
 INV_X1 _20985_ (.A(_15161_),
    .ZN(_15801_));
 INV_X1 _20986_ (.A(_15152_),
    .ZN(_15200_));
 INV_X1 _20987_ (.A(_15172_),
    .ZN(_15802_));
 INV_X1 _20988_ (.A(_15238_),
    .ZN(_15806_));
 INV_X1 _20989_ (.A(_15249_),
    .ZN(_15808_));
 INV_X1 _20990_ (.A(_15254_),
    .ZN(_15255_));
 INV_X1 _20991_ (.A(_15261_),
    .ZN(_15265_));
 INV_X1 _20992_ (.A(_15278_),
    .ZN(_15812_));
 INV_X1 _20993_ (.A(_15228_),
    .ZN(_15279_));
 INV_X1 _20994_ (.A(_15289_),
    .ZN(_15814_));
 INV_X1 _20995_ (.A(_15293_),
    .ZN(_15294_));
 INV_X1 _20996_ (.A(_15324_),
    .ZN(_15820_));
 INV_X1 _20997_ (.A(_15351_),
    .ZN(_15827_));
 INV_X1 _20998_ (.A(_15928_),
    .ZN(_15924_));
 INV_X1 _20999_ (.A(_15944_),
    .ZN(_15940_));
 INV_X2 _21000_ (.A(_15992_),
    .ZN(_15988_));
 INV_X1 _21001_ (.A(_16000_),
    .ZN(_15996_));
 INV_X1 _21002_ (.A(_16008_),
    .ZN(_16004_));
 INV_X1 _21003_ (.A(_16016_),
    .ZN(_16012_));
 INV_X1 _21004_ (.A(_16032_),
    .ZN(_16028_));
 INV_X1 _21005_ (.A(_16040_),
    .ZN(_16036_));
 INV_X1 _21006_ (.A(_16048_),
    .ZN(_16044_));
 INV_X1 _21007_ (.A(_16080_),
    .ZN(_16076_));
 BUF_X4 _21008_ (.A(_03620_),
    .Z(_04153_));
 BUF_X4 _21009_ (.A(_04153_),
    .Z(_16084_));
 BUF_X4 _21010_ (.A(_03957_),
    .Z(_04154_));
 BUF_X2 _21011_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Z(_04155_));
 BUF_X4 _21012_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_04156_));
 BUF_X4 _21013_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_04157_));
 BUF_X4 _21014_ (.A(_04157_),
    .Z(_04158_));
 OAI221_X2 _21015_ (.A(_04154_),
    .B1(_04155_),
    .B2(_04156_),
    .C1(_04158_),
    .C2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_04159_));
 NOR2_X2 _21016_ (.A1(_11420_),
    .A2(_11422_),
    .ZN(_04160_));
 OAI22_X2 _21017_ (.A1(_11422_),
    .A2(_11424_),
    .B1(_03877_),
    .B2(_04160_),
    .ZN(_04161_));
 NAND3_X2 _21018_ (.A1(_00134_),
    .A2(_04159_),
    .A3(_04161_),
    .ZN(_04162_));
 INV_X1 _21019_ (.A(_04162_),
    .ZN(_04163_));
 NAND2_X4 _21020_ (.A1(_00133_),
    .A2(_04163_),
    .ZN(_04164_));
 INV_X2 _21021_ (.A(_04164_),
    .ZN(_16107_));
 OR3_X1 _21022_ (.A1(_00185_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04165_));
 OAI21_X1 _21023_ (.A(_04165_),
    .B1(_04043_),
    .B2(_15849_),
    .ZN(_15370_));
 OR3_X1 _21024_ (.A1(_00217_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04166_));
 OAI21_X2 _21025_ (.A(_04166_),
    .B1(_04043_),
    .B2(_15838_),
    .ZN(_14066_));
 OR3_X1 _21026_ (.A1(_00556_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04167_));
 OAI21_X1 _21027_ (.A(_04167_),
    .B1(_15856_),
    .B2(_04090_),
    .ZN(_15376_));
 OR3_X1 _21028_ (.A1(_00557_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04168_));
 OAI21_X1 _21029_ (.A(_04168_),
    .B1(_15861_),
    .B2(_04090_),
    .ZN(_15380_));
 OR3_X1 _21030_ (.A1(_00558_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04169_));
 OAI21_X1 _21031_ (.A(_04169_),
    .B1(_15872_),
    .B2(_04090_),
    .ZN(_15384_));
 OR3_X1 _21032_ (.A1(_00559_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04170_));
 BUF_X2 _21033_ (.A(_04028_),
    .Z(_04171_));
 OAI21_X1 _21034_ (.A(_04170_),
    .B1(_15881_),
    .B2(_04171_),
    .ZN(_15388_));
 OR3_X1 _21035_ (.A1(_00560_),
    .A2(_04134_),
    .A3(_04135_),
    .ZN(_04172_));
 OAI21_X1 _21036_ (.A(_04172_),
    .B1(_15889_),
    .B2(_04171_),
    .ZN(_15392_));
 XNOR2_X1 _21037_ (.A(_15896_),
    .B(_04030_),
    .ZN(_04173_));
 OAI222_X2 _21038_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .B2(_04033_),
    .C1(_03723_),
    .C2(_03402_),
    .ZN(_04174_));
 NOR2_X1 _21039_ (.A1(_04071_),
    .A2(_04174_),
    .ZN(_04175_));
 AOI21_X1 _21040_ (.A(_04175_),
    .B1(_04071_),
    .B2(_11202_),
    .ZN(_04176_));
 MUX2_X1 _21041_ (.A(_04173_),
    .B(_04176_),
    .S(_04132_),
    .Z(_15396_));
 CLKBUF_X2 _21042_ (.A(_11409_),
    .Z(_04177_));
 CLKBUF_X2 _21043_ (.A(_04107_),
    .Z(_04178_));
 OR3_X1 _21044_ (.A1(_00562_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04179_));
 OAI21_X1 _21045_ (.A(_04179_),
    .B1(_15905_),
    .B2(_04171_),
    .ZN(_15400_));
 OR3_X1 _21046_ (.A1(_00563_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04180_));
 OAI21_X1 _21047_ (.A(_04180_),
    .B1(_15913_),
    .B2(_04171_),
    .ZN(_15404_));
 OR3_X1 _21048_ (.A1(_00564_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04181_));
 OAI21_X1 _21049_ (.A(_04181_),
    .B1(_15921_),
    .B2(_04171_),
    .ZN(_15408_));
 XNOR2_X1 _21050_ (.A(_15929_),
    .B(_04030_),
    .ZN(_04182_));
 OAI222_X2 _21051_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .B2(_04033_),
    .C1(_11398_),
    .C2(_04055_),
    .ZN(_04183_));
 MUX2_X1 _21052_ (.A(_03743_),
    .B(_04183_),
    .S(_03406_),
    .Z(_04184_));
 MUX2_X1 _21053_ (.A(_04182_),
    .B(_04184_),
    .S(_04132_),
    .Z(_15412_));
 XNOR2_X1 _21054_ (.A(_04050_),
    .B(_15937_),
    .ZN(_04185_));
 OAI222_X2 _21055_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .B2(_04054_),
    .C1(_10868_),
    .C2(_04112_),
    .ZN(_04186_));
 NAND2_X1 _21056_ (.A1(_04128_),
    .A2(_04186_),
    .ZN(_04187_));
 OAI21_X1 _21057_ (.A(_04187_),
    .B1(_04141_),
    .B2(_11993_),
    .ZN(_04188_));
 MUX2_X1 _21058_ (.A(_04185_),
    .B(_04188_),
    .S(_04132_),
    .Z(_15416_));
 XNOR2_X1 _21059_ (.A(_04050_),
    .B(_15945_),
    .ZN(_04189_));
 OAI222_X2 _21060_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .B2(_04054_),
    .C1(_12075_),
    .C2(_04112_),
    .ZN(_04190_));
 NAND2_X1 _21061_ (.A1(_04128_),
    .A2(_04190_),
    .ZN(_04191_));
 OAI21_X1 _21062_ (.A(_04191_),
    .B1(_04141_),
    .B2(_12044_),
    .ZN(_04192_));
 MUX2_X1 _21063_ (.A(_04189_),
    .B(_04192_),
    .S(_04132_),
    .Z(_15420_));
 OR3_X1 _21064_ (.A1(_04026_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04193_));
 OAI21_X1 _21065_ (.A(_04193_),
    .B1(_15952_),
    .B2(_04171_),
    .ZN(_15424_));
 OR3_X1 _21066_ (.A1(_00659_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04194_));
 OAI21_X1 _21067_ (.A(_04194_),
    .B1(_15957_),
    .B2(_04171_),
    .ZN(_15428_));
 OR3_X1 _21068_ (.A1(_03670_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04195_));
 OAI21_X1 _21069_ (.A(_04195_),
    .B1(_15968_),
    .B2(_04171_),
    .ZN(_15432_));
 OR3_X1 _21070_ (.A1(_03800_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04196_));
 OAI21_X1 _21071_ (.A(_04196_),
    .B1(_15976_),
    .B2(_04171_),
    .ZN(_15436_));
 OR3_X1 _21072_ (.A1(_03804_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04197_));
 OAI21_X1 _21073_ (.A(_04197_),
    .B1(_15981_),
    .B2(_04171_),
    .ZN(_15440_));
 XNOR2_X1 _21074_ (.A(net317),
    .B(_15993_),
    .ZN(_04198_));
 OAI222_X2 _21075_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .B2(_04054_),
    .C1(_12589_),
    .C2(_04112_),
    .ZN(_04199_));
 NAND2_X1 _21076_ (.A1(_04128_),
    .A2(_04199_),
    .ZN(_04200_));
 OAI21_X1 _21077_ (.A(_04200_),
    .B1(_04141_),
    .B2(net349),
    .ZN(_04201_));
 MUX2_X1 _21078_ (.A(_04198_),
    .B(_04201_),
    .S(_04132_),
    .Z(_15444_));
 OR3_X1 _21079_ (.A1(_03808_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04202_));
 OAI21_X1 _21080_ (.A(_04202_),
    .B1(_15997_),
    .B2(_04029_),
    .ZN(_15448_));
 XNOR2_X1 _21081_ (.A(_04117_),
    .B(_16008_),
    .ZN(_04203_));
 OAI222_X2 _21082_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .B2(_04054_),
    .C1(net361),
    .C2(_04055_),
    .ZN(_04204_));
 NAND2_X1 _21083_ (.A1(_04128_),
    .A2(_04204_),
    .ZN(_04205_));
 OAI21_X1 _21084_ (.A(_04205_),
    .B1(_04141_),
    .B2(_12725_),
    .ZN(_04206_));
 MUX2_X1 _21085_ (.A(_04203_),
    .B(_04206_),
    .S(_04132_),
    .Z(_15452_));
 OR3_X1 _21086_ (.A1(_03813_),
    .A2(_04177_),
    .A3(_04178_),
    .ZN(_04207_));
 OAI21_X1 _21087_ (.A(_04207_),
    .B1(_16013_),
    .B2(_04029_),
    .ZN(_15456_));
 OR3_X1 _21088_ (.A1(_03815_),
    .A2(_11409_),
    .A3(_04034_),
    .ZN(_04208_));
 OAI21_X1 _21089_ (.A(_04208_),
    .B1(_16024_),
    .B2(_04029_),
    .ZN(_15460_));
 XNOR2_X1 _21090_ (.A(_04117_),
    .B(_16032_),
    .ZN(_04209_));
 OAI222_X2 _21091_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .B2(_04054_),
    .C1(_03733_),
    .C2(_04055_),
    .ZN(_04210_));
 NAND2_X1 _21092_ (.A1(_04128_),
    .A2(_04210_),
    .ZN(_04211_));
 OAI21_X1 _21093_ (.A(_04211_),
    .B1(_04141_),
    .B2(_12985_),
    .ZN(_04212_));
 MUX2_X1 _21094_ (.A(_04209_),
    .B(_04212_),
    .S(_04028_),
    .Z(_15464_));
 XNOR2_X1 _21095_ (.A(_04117_),
    .B(_16037_),
    .ZN(_04213_));
 OAI222_X2 _21096_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .B2(_04054_),
    .C1(_13097_),
    .C2(_04055_),
    .ZN(_04214_));
 NAND2_X1 _21097_ (.A1(_04128_),
    .A2(_04214_),
    .ZN(_04215_));
 OAI21_X1 _21098_ (.A(_04215_),
    .B1(_04141_),
    .B2(_13061_),
    .ZN(_04216_));
 MUX2_X1 _21099_ (.A(_04213_),
    .B(_04216_),
    .S(_04028_),
    .Z(_15468_));
 OR3_X1 _21100_ (.A1(_01000_),
    .A2(_11409_),
    .A3(_04034_),
    .ZN(_04217_));
 OAI21_X2 _21101_ (.A(_04217_),
    .B1(_16045_),
    .B2(_04029_),
    .ZN(_15472_));
 OR3_X1 _21102_ (.A1(_03824_),
    .A2(_11409_),
    .A3(_04034_),
    .ZN(_04218_));
 OAI21_X2 _21103_ (.A(_04218_),
    .B1(_16056_),
    .B2(_04029_),
    .ZN(_15476_));
 XNOR2_X1 _21104_ (.A(_04117_),
    .B(_16061_),
    .ZN(_04219_));
 OAI222_X2 _21105_ (.A1(_04138_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .B2(_04054_),
    .C1(_03762_),
    .C2(_04055_),
    .ZN(_04220_));
 NAND2_X1 _21106_ (.A1(_04040_),
    .A2(_04220_),
    .ZN(_04221_));
 OAI21_X1 _21107_ (.A(_04221_),
    .B1(_04141_),
    .B2(_13314_),
    .ZN(_04222_));
 MUX2_X1 _21108_ (.A(_04219_),
    .B(_04222_),
    .S(_04028_),
    .Z(_15480_));
 OR3_X1 _21109_ (.A1(_01093_),
    .A2(_11409_),
    .A3(_04034_),
    .ZN(_04223_));
 OAI21_X2 _21110_ (.A(_04223_),
    .B1(_16072_),
    .B2(_04029_),
    .ZN(_15484_));
 XNOR2_X1 _21111_ (.A(_11863_),
    .B(_16077_),
    .ZN(_04224_));
 OAI222_X2 _21112_ (.A1(_04044_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .B2(_04054_),
    .C1(_03311_),
    .C2(_04055_),
    .ZN(_04225_));
 NAND2_X1 _21113_ (.A1(_04040_),
    .A2(_04225_),
    .ZN(_04226_));
 OAI21_X1 _21114_ (.A(_04226_),
    .B1(_04035_),
    .B2(_03275_),
    .ZN(_04227_));
 MUX2_X1 _21115_ (.A(_04224_),
    .B(_04227_),
    .S(_04028_),
    .Z(_15488_));
 INV_X1 _21116_ (.A(_15526_),
    .ZN(_15523_));
 INV_X1 _21117_ (.A(_14073_),
    .ZN(_15554_));
 INV_X1 _21118_ (.A(_14072_),
    .ZN(_15558_));
 INV_X1 _21119_ (.A(_14083_),
    .ZN(_15570_));
 INV_X1 _21120_ (.A(_14077_),
    .ZN(_15569_));
 INV_X1 _21121_ (.A(_14093_),
    .ZN(_14095_));
 INV_X1 _21122_ (.A(_14082_),
    .ZN(_14096_));
 INV_X1 _21123_ (.A(_14103_),
    .ZN(_15587_));
 INV_X1 _21124_ (.A(_14102_),
    .ZN(_14123_));
 INV_X1 _21125_ (.A(_14120_),
    .ZN(_15617_));
 INV_X1 _21126_ (.A(_14149_),
    .ZN(_14156_));
 INV_X1 _21127_ (.A(_14138_),
    .ZN(_15623_));
 INV_X1 _21128_ (.A(_14143_),
    .ZN(_15629_));
 INV_X1 _21129_ (.A(_14165_),
    .ZN(_15638_));
 INV_X1 _21130_ (.A(_14170_),
    .ZN(_14205_));
 INV_X1 _21131_ (.A(_14175_),
    .ZN(_15642_));
 INV_X1 _21132_ (.A(_14188_),
    .ZN(_15650_));
 INV_X1 _21133_ (.A(_14201_),
    .ZN(_14240_));
 INV_X1 _21134_ (.A(_14219_),
    .ZN(_15663_));
 INV_X1 _21135_ (.A(_14282_),
    .ZN(_15670_));
 INV_X1 _21136_ (.A(_14246_),
    .ZN(_15674_));
 INV_X2 _21137_ (.A(_14325_),
    .ZN(_15684_));
 INV_X1 _21138_ (.A(_14286_),
    .ZN(_15692_));
 INV_X1 _21139_ (.A(_14310_),
    .ZN(_15696_));
 INV_X1 _21140_ (.A(_14302_),
    .ZN(_14361_));
 INV_X1 _21141_ (.A(_14324_),
    .ZN(_15698_));
 INV_X1 _21142_ (.A(_14384_),
    .ZN(_15701_));
 INV_X1 _21143_ (.A(_14358_),
    .ZN(_15703_));
 INV_X1 _21144_ (.A(_14345_),
    .ZN(_14415_));
 INV_X1 _21145_ (.A(_14370_),
    .ZN(_15705_));
 INV_X1 _21146_ (.A(_14432_),
    .ZN(_15709_));
 INV_X2 _21147_ (.A(_14455_),
    .ZN(_14457_));
 INV_X1 _21148_ (.A(_14412_),
    .ZN(_15713_));
 INV_X1 _21149_ (.A(_14399_),
    .ZN(_14470_));
 INV_X1 _21150_ (.A(_14426_),
    .ZN(_15715_));
 INV_X2 _21151_ (.A(_14513_),
    .ZN(_14515_));
 INV_X1 _21152_ (.A(_14467_),
    .ZN(_15722_));
 INV_X1 _21153_ (.A(_14454_),
    .ZN(_14527_));
 INV_X1 _21154_ (.A(_14480_),
    .ZN(_15724_));
 INV_X1 _21155_ (.A(_14524_),
    .ZN(_14595_));
 INV_X1 _21156_ (.A(_14537_),
    .ZN(_15728_));
 INV_X1 _21157_ (.A(_14591_),
    .ZN(_15734_));
 INV_X1 _21158_ (.A(_14607_),
    .ZN(_15737_));
 INV_X1 _21159_ (.A(_14658_),
    .ZN(_15741_));
 INV_X1 _21160_ (.A(_14667_),
    .ZN(_15743_));
 INV_X1 _21161_ (.A(_14715_),
    .ZN(_15747_));
 INV_X1 _21162_ (.A(_14705_),
    .ZN(_14775_));
 INV_X1 _21163_ (.A(_14725_),
    .ZN(_15749_));
 INV_X1 _21164_ (.A(_14841_),
    .ZN(_15755_));
 INV_X1 _21165_ (.A(_14829_),
    .ZN(_15759_));
 INV_X1 _21166_ (.A(_14820_),
    .ZN(_14885_));
 INV_X1 _21167_ (.A(_14840_),
    .ZN(_15761_));
 INV_X1 _21168_ (.A(_14921_),
    .ZN(_14923_));
 INV_X1 _21169_ (.A(_14948_),
    .ZN(_15767_));
 INV_X1 _21170_ (.A(_14936_),
    .ZN(_15771_));
 INV_X1 _21171_ (.A(_14947_),
    .ZN(_15773_));
 INV_X1 _21172_ (.A(_14980_),
    .ZN(_15039_));
 INV_X1 _21173_ (.A(_15047_),
    .ZN(_15779_));
 INV_X1 _21174_ (.A(_15079_),
    .ZN(_15783_));
 INV_X1 _21175_ (.A(_15046_),
    .ZN(_15785_));
 INV_X1 _21176_ (.A(_15078_),
    .ZN(_15789_));
 INV_X1 _21177_ (.A(_15089_),
    .ZN(_15791_));
 INV_X1 _21178_ (.A(_15173_),
    .ZN(_15797_));
 INV_X1 _21179_ (.A(_15210_),
    .ZN(_15803_));
 INV_X1 _21180_ (.A(_15198_),
    .ZN(_15807_));
 INV_X1 _21181_ (.A(_15189_),
    .ZN(_15240_));
 INV_X1 _21182_ (.A(_15209_),
    .ZN(_15809_));
 INV_X1 _21183_ (.A(_15214_),
    .ZN(_15256_));
 INV_X1 _21184_ (.A(_15224_),
    .ZN(_15266_));
 INV_X1 _21185_ (.A(_15237_),
    .ZN(_15813_));
 INV_X1 _21186_ (.A(_15248_),
    .ZN(_15815_));
 INV_X1 _21187_ (.A(_15253_),
    .ZN(_15295_));
 INV_X1 _21188_ (.A(_15260_),
    .ZN(_15302_));
 INV_X1 _21189_ (.A(_15314_),
    .ZN(_15819_));
 INV_X1 _21190_ (.A(_15277_),
    .ZN(_15818_));
 INV_X1 _21191_ (.A(_15288_),
    .ZN(_15821_));
 INV_X1 _21192_ (.A(_15292_),
    .ZN(_15329_));
 INV_X1 _21193_ (.A(_15313_),
    .ZN(_15825_));
 INV_X1 _21194_ (.A(_15323_),
    .ZN(_15828_));
 INV_X1 _21195_ (.A(_15881_),
    .ZN(_15877_));
 INV_X1 _21196_ (.A(_15889_),
    .ZN(_15885_));
 INV_X1 _21197_ (.A(_16021_),
    .ZN(_16025_));
 INV_X1 _21198_ (.A(_16037_),
    .ZN(_16041_));
 INV_X2 _21199_ (.A(_16045_),
    .ZN(_16049_));
 INV_X1 _21200_ (.A(_16053_),
    .ZN(_16057_));
 INV_X1 _21201_ (.A(_16061_),
    .ZN(_16065_));
 INV_X1 _21202_ (.A(_16069_),
    .ZN(_16073_));
 INV_X1 _21203_ (.A(_16077_),
    .ZN(_16081_));
 INV_X1 _21204_ (.A(_15586_),
    .ZN(_14100_));
 INV_X1 _21205_ (.A(_15598_),
    .ZN(_14118_));
 INV_X1 _21206_ (.A(_15615_),
    .ZN(_14140_));
 INV_X1 _21207_ (.A(_15625_),
    .ZN(_14167_));
 INV_X1 _21208_ (.A(_15627_),
    .ZN(_14173_));
 INV_X1 _21209_ (.A(_15640_),
    .ZN(_14198_));
 INV_X1 _21210_ (.A(_15656_),
    .ZN(_14231_));
 INV_X1 _21211_ (.A(_15669_),
    .ZN(_14271_));
 INV_X1 _21212_ (.A(_15682_),
    .ZN(_14314_));
 INV_X1 _21213_ (.A(_15735_),
    .ZN(_14660_));
 INV_X1 _21214_ (.A(_15660_),
    .ZN(_14301_));
 INV_X1 _21215_ (.A(_15675_),
    .ZN(_14344_));
 INV_X1 _21216_ (.A(_15689_),
    .ZN(_14382_));
 INV_X1 _21217_ (.A(_15693_),
    .ZN(_14398_));
 NOR3_X1 _21218_ (.A1(_11430_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .A3(_11406_),
    .ZN(_04228_));
 AND2_X4 _21219_ (.A1(_11403_),
    .A2(_04228_),
    .ZN(_04229_));
 OAI33_X1 _21220_ (.A1(_10341_),
    .A2(_10372_),
    .A3(_10299_),
    .B1(_10333_),
    .B2(_10384_),
    .B3(_10364_),
    .ZN(_04230_));
 AOI21_X4 _21221_ (.A(_03493_),
    .B1(_04230_),
    .B2(_10312_),
    .ZN(_04231_));
 NOR2_X2 _21222_ (.A1(_04229_),
    .A2(_04231_),
    .ZN(_04232_));
 AND3_X1 _21223_ (.A1(_10921_),
    .A2(_03533_),
    .A3(_03514_),
    .ZN(_04233_));
 OAI21_X1 _21224_ (.A(_03527_),
    .B1(_11071_),
    .B2(_10920_),
    .ZN(_04234_));
 OAI221_X2 _21225_ (.A(_04233_),
    .B1(_04234_),
    .B2(_15869_),
    .C1(_03506_),
    .C2(_03505_),
    .ZN(_04235_));
 NAND2_X2 _21226_ (.A1(_03554_),
    .A2(_03533_),
    .ZN(_04236_));
 OAI21_X2 _21227_ (.A(_04235_),
    .B1(_03551_),
    .B2(_04236_),
    .ZN(_04237_));
 OAI211_X4 _21228_ (.A(_10921_),
    .B(_03491_),
    .C1(_11352_),
    .C2(_11321_),
    .ZN(_04238_));
 NOR2_X2 _21229_ (.A1(_15916_),
    .A2(_04238_),
    .ZN(_04239_));
 OAI21_X1 _21230_ (.A(_04239_),
    .B1(_03558_),
    .B2(_03561_),
    .ZN(_04240_));
 NAND3_X1 _21231_ (.A1(_03537_),
    .A2(_04239_),
    .A3(_03569_),
    .ZN(_04241_));
 NAND2_X1 _21232_ (.A1(_04240_),
    .A2(_04241_),
    .ZN(_04242_));
 NAND2_X1 _21233_ (.A1(_15884_),
    .A2(_15896_),
    .ZN(_04243_));
 OR4_X4 _21234_ (.A1(_15916_),
    .A2(_04238_),
    .A3(_03524_),
    .A4(_04243_),
    .ZN(_04244_));
 OAI21_X2 _21235_ (.A(_03506_),
    .B1(_03530_),
    .B2(_03499_),
    .ZN(_04245_));
 AOI21_X2 _21236_ (.A(_04244_),
    .B1(_04245_),
    .B2(_03575_),
    .ZN(_04246_));
 OAI21_X4 _21237_ (.A(_04239_),
    .B1(_03584_),
    .B2(_03582_),
    .ZN(_04247_));
 NOR2_X2 _21238_ (.A1(_10919_),
    .A2(_15884_),
    .ZN(_04248_));
 AND4_X2 _21239_ (.A1(_15929_),
    .A2(_03491_),
    .A3(_04248_),
    .A4(_03587_),
    .ZN(_04249_));
 NOR3_X1 _21240_ (.A1(_10919_),
    .A2(_15880_),
    .A3(_03555_),
    .ZN(_04250_));
 OAI211_X2 _21241_ (.A(_04249_),
    .B(_04250_),
    .C1(_03506_),
    .C2(_03580_),
    .ZN(_04251_));
 AOI21_X1 _21242_ (.A(_04238_),
    .B1(_15916_),
    .B2(_11065_),
    .ZN(_04252_));
 NAND4_X1 _21243_ (.A1(_03530_),
    .A2(_03554_),
    .A3(_03556_),
    .A4(_04252_),
    .ZN(_04253_));
 AND2_X1 _21244_ (.A1(_04251_),
    .A2(_04253_),
    .ZN(_04254_));
 NOR4_X4 _21245_ (.A1(_10934_),
    .A2(_10975_),
    .A3(_15864_),
    .A4(_03596_),
    .ZN(_04255_));
 NAND3_X2 _21246_ (.A1(_03514_),
    .A2(_04255_),
    .A3(_03595_),
    .ZN(_04256_));
 NAND3_X1 _21247_ (.A1(_15884_),
    .A2(_03542_),
    .A3(_03599_),
    .ZN(_04257_));
 OR4_X1 _21248_ (.A1(_15920_),
    .A2(_04238_),
    .A3(_03580_),
    .A4(_04257_),
    .ZN(_04258_));
 NAND4_X2 _21249_ (.A1(_04247_),
    .A2(_04254_),
    .A3(_04256_),
    .A4(_04258_),
    .ZN(_04259_));
 NOR4_X4 _21250_ (.A1(_04237_),
    .A2(_04242_),
    .A3(_04246_),
    .A4(_04259_),
    .ZN(_04260_));
 OAI21_X4 _21251_ (.A(_10922_),
    .B1(_03508_),
    .B2(_04260_),
    .ZN(_04261_));
 AND3_X1 _21252_ (.A1(_03439_),
    .A2(_04232_),
    .A3(_04261_),
    .ZN(_04262_));
 BUF_X4 _21253_ (.A(_04262_),
    .Z(_04263_));
 BUF_X4 _21254_ (.A(_11482_),
    .Z(_04264_));
 NAND2_X4 _21255_ (.A1(_11512_),
    .A2(_11918_),
    .ZN(_04265_));
 NAND2_X2 _21256_ (.A1(_11492_),
    .A2(_11508_),
    .ZN(_04266_));
 NOR2_X4 _21257_ (.A1(_11510_),
    .A2(_04266_),
    .ZN(_04267_));
 INV_X1 _21258_ (.A(_11505_),
    .ZN(_04268_));
 NAND2_X2 _21259_ (.A1(_11476_),
    .A2(_04268_),
    .ZN(_04269_));
 AOI21_X4 _21260_ (.A(net301),
    .B1(_04267_),
    .B2(_04269_),
    .ZN(_04270_));
 CLKBUF_X3 _21261_ (.A(_15359_),
    .Z(_04271_));
 INV_X1 _21262_ (.A(_04271_),
    .ZN(_04272_));
 BUF_X4 _21263_ (.A(_11500_),
    .Z(_04273_));
 NOR2_X2 _21264_ (.A1(_04272_),
    .A2(_04273_),
    .ZN(_04274_));
 NOR4_X4 _21265_ (.A1(_04264_),
    .A2(_04265_),
    .A3(_04270_),
    .A4(_04274_),
    .ZN(_04275_));
 BUF_X4 _21266_ (.A(_04275_),
    .Z(_04276_));
 INV_X1 _21267_ (.A(_15836_),
    .ZN(_04277_));
 AOI211_X2 _21268_ (.A(_04277_),
    .B(_15864_),
    .C1(_11067_),
    .C2(_11070_),
    .ZN(_04278_));
 OAI21_X4 _21269_ (.A(_15873_),
    .B1(_04278_),
    .B2(_10333_),
    .ZN(_04279_));
 OR3_X4 _21270_ (.A1(_10333_),
    .A2(_11065_),
    .A3(_04278_),
    .ZN(_04280_));
 AND2_X2 _21271_ (.A1(_04279_),
    .A2(_04280_),
    .ZN(_04281_));
 BUF_X4 _21272_ (.A(_04281_),
    .Z(_04282_));
 AOI21_X2 _21273_ (.A(_10737_),
    .B1(_10476_),
    .B2(_10396_),
    .ZN(_04283_));
 AOI22_X4 _21274_ (.A1(_10333_),
    .A2(_15860_),
    .B1(_11071_),
    .B2(_04283_),
    .ZN(_04284_));
 OAI21_X2 _21275_ (.A(_10673_),
    .B1(_10317_),
    .B2(net345),
    .ZN(_04285_));
 AND2_X1 _21276_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_10354_),
    .ZN(_04286_));
 MUX2_X1 _21277_ (.A(net357),
    .B(_04286_),
    .S(_10376_),
    .Z(_04287_));
 AOI221_X2 _21278_ (.A(_10403_),
    .B1(_10389_),
    .B2(_04287_),
    .C1(_10932_),
    .C2(_10394_),
    .ZN(_04288_));
 OAI21_X2 _21279_ (.A(_10736_),
    .B1(_04285_),
    .B2(_04288_),
    .ZN(_04289_));
 OAI221_X2 _21280_ (.A(_15864_),
    .B1(_04289_),
    .B2(_15853_),
    .C1(_10306_),
    .C2(_10305_),
    .ZN(_04290_));
 AND2_X1 _21281_ (.A1(_04284_),
    .A2(_04290_),
    .ZN(_04291_));
 CLKBUF_X3 _21282_ (.A(_04291_),
    .Z(_04292_));
 CLKBUF_X3 _21283_ (.A(_04292_),
    .Z(_04293_));
 NAND2_X2 _21284_ (.A1(_15837_),
    .A2(_10368_),
    .ZN(_04294_));
 CLKBUF_X3 _21285_ (.A(_04294_),
    .Z(_04295_));
 AOI22_X4 _21286_ (.A1(_04277_),
    .A2(_10368_),
    .B1(_11070_),
    .B2(_11067_),
    .ZN(_04296_));
 NOR4_X4 _21287_ (.A1(_15836_),
    .A2(_10333_),
    .A3(_10934_),
    .A4(_10975_),
    .ZN(_04297_));
 OAI221_X2 _21288_ (.A(_04295_),
    .B1(_04296_),
    .B2(_04297_),
    .C1(_10368_),
    .C2(_15834_),
    .ZN(_04298_));
 AOI21_X2 _21289_ (.A(_04282_),
    .B1(_04293_),
    .B2(_04298_),
    .ZN(_04299_));
 INV_X4 _21290_ (.A(_04264_),
    .ZN(_04300_));
 NOR3_X4 _21291_ (.A1(_11510_),
    .A2(_11862_),
    .A3(_04266_),
    .ZN(_04301_));
 NAND3_X4 _21292_ (.A1(_04271_),
    .A2(_04300_),
    .A3(_04301_),
    .ZN(_04302_));
 MUX2_X2 _21293_ (.A(_15842_),
    .B(_15496_),
    .S(_04302_),
    .Z(_04303_));
 NAND2_X2 _21294_ (.A1(_11486_),
    .A2(_04300_),
    .ZN(_04304_));
 NOR3_X2 _21295_ (.A1(_04273_),
    .A2(_04304_),
    .A3(_04265_),
    .ZN(_04305_));
 AND2_X2 _21296_ (.A1(_04303_),
    .A2(_04305_),
    .ZN(_04306_));
 BUF_X4 _21297_ (.A(_04306_),
    .Z(_04307_));
 CLKBUF_X3 _21298_ (.A(_04282_),
    .Z(_04308_));
 NOR3_X1 _21299_ (.A1(_15835_),
    .A2(_04297_),
    .A3(_04296_),
    .ZN(_04309_));
 OR3_X2 _21300_ (.A1(_04272_),
    .A2(_11482_),
    .A3(_11484_),
    .ZN(_04310_));
 OR2_X1 _21301_ (.A1(_11500_),
    .A2(_04310_),
    .ZN(_04311_));
 BUF_X4 _21302_ (.A(_04311_),
    .Z(_04312_));
 BUF_X4 _21303_ (.A(_04312_),
    .Z(_04313_));
 MUX2_X1 _21304_ (.A(_15856_),
    .B(_16072_),
    .S(_04313_),
    .Z(_04314_));
 NAND3_X2 _21305_ (.A1(_10333_),
    .A2(_10396_),
    .A3(_10476_),
    .ZN(_04315_));
 BUF_X2 _21306_ (.A(_04315_),
    .Z(_04316_));
 AOI21_X2 _21307_ (.A(_04314_),
    .B1(_04295_),
    .B2(_04316_),
    .ZN(_04317_));
 NOR3_X4 _21308_ (.A1(_10368_),
    .A2(_04288_),
    .A3(_04285_),
    .ZN(_04318_));
 AND2_X1 _21309_ (.A1(_15837_),
    .A2(_10368_),
    .ZN(_04319_));
 CLKBUF_X3 _21310_ (.A(_04319_),
    .Z(_04320_));
 MUX2_X1 _21311_ (.A(_15872_),
    .B(_16056_),
    .S(_04313_),
    .Z(_04321_));
 NOR3_X1 _21312_ (.A1(_04318_),
    .A2(_04320_),
    .A3(_04321_),
    .ZN(_04322_));
 OAI21_X1 _21313_ (.A(_04309_),
    .B1(_04317_),
    .B2(_04322_),
    .ZN(_04323_));
 MUX2_X1 _21314_ (.A(_15905_),
    .B(_16024_),
    .S(_04312_),
    .Z(_04324_));
 MUX2_X1 _21315_ (.A(_15913_),
    .B(_16013_),
    .S(_04312_),
    .Z(_04325_));
 MUX2_X1 _21316_ (.A(_04324_),
    .B(_04325_),
    .S(_10736_),
    .Z(_04326_));
 MUX2_X1 _21317_ (.A(_15889_),
    .B(_16040_),
    .S(_04312_),
    .Z(_04327_));
 MUX2_X1 _21318_ (.A(_15897_),
    .B(_16029_),
    .S(_04312_),
    .Z(_04328_));
 MUX2_X1 _21319_ (.A(_04327_),
    .B(_04328_),
    .S(_10736_),
    .Z(_04329_));
 NAND2_X4 _21320_ (.A1(_04315_),
    .A2(_04294_),
    .ZN(_04330_));
 MUX2_X1 _21321_ (.A(_04326_),
    .B(_04329_),
    .S(_04330_),
    .Z(_04331_));
 NOR2_X4 _21322_ (.A1(_04297_),
    .A2(_04296_),
    .ZN(_04332_));
 BUF_X4 _21323_ (.A(_04332_),
    .Z(_04333_));
 MUX2_X1 _21324_ (.A(_15881_),
    .B(_16045_),
    .S(_04313_),
    .Z(_04334_));
 NOR3_X1 _21325_ (.A1(_04318_),
    .A2(_04320_),
    .A3(_04334_),
    .ZN(_04335_));
 MUX2_X1 _21326_ (.A(_15861_),
    .B(_16064_),
    .S(_04302_),
    .Z(_04336_));
 AOI21_X1 _21327_ (.A(_04336_),
    .B1(_04294_),
    .B2(_04315_),
    .ZN(_04337_));
 NOR2_X1 _21328_ (.A1(_04335_),
    .A2(_04337_),
    .ZN(_04338_));
 NAND2_X1 _21329_ (.A1(_15835_),
    .A2(_04333_),
    .ZN(_04339_));
 OAI221_X2 _21330_ (.A(_04323_),
    .B1(_04331_),
    .B2(_04333_),
    .C1(_04338_),
    .C2(_04339_),
    .ZN(_04340_));
 NOR2_X1 _21331_ (.A1(_15845_),
    .A2(_04313_),
    .ZN(_04341_));
 BUF_X4 _21332_ (.A(_04313_),
    .Z(_04342_));
 AOI21_X2 _21333_ (.A(_04341_),
    .B1(_04342_),
    .B2(_16080_),
    .ZN(_04343_));
 MUX2_X1 _21334_ (.A(_04303_),
    .B(_04343_),
    .S(_10739_),
    .Z(_04344_));
 OR2_X1 _21335_ (.A1(_04298_),
    .A2(_04344_),
    .ZN(_04345_));
 MUX2_X1 _21336_ (.A(_04340_),
    .B(_04345_),
    .S(_04293_),
    .Z(_04346_));
 OAI221_X2 _21337_ (.A(_04276_),
    .B1(_04299_),
    .B2(_04307_),
    .C1(_04308_),
    .C2(_04346_),
    .ZN(_04347_));
 NOR2_X2 _21338_ (.A1(_04300_),
    .A2(_04265_),
    .ZN(_04348_));
 MUX2_X1 _21339_ (.A(net297),
    .B(_04271_),
    .S(_04273_),
    .Z(_04349_));
 AND2_X2 _21340_ (.A1(_04348_),
    .A2(_04349_),
    .ZN(_04350_));
 BUF_X4 _21341_ (.A(_04350_),
    .Z(_04351_));
 CLKBUF_X3 _21342_ (.A(_04351_),
    .Z(_04352_));
 CLKBUF_X3 _21343_ (.A(_04352_),
    .Z(_04353_));
 NAND3_X4 _21344_ (.A1(_04264_),
    .A2(_11512_),
    .A3(_11918_),
    .ZN(_04354_));
 NAND2_X1 _21345_ (.A1(_04271_),
    .A2(_04267_),
    .ZN(_04355_));
 NOR2_X2 _21346_ (.A1(net297),
    .A2(net301),
    .ZN(_04356_));
 NAND3_X2 _21347_ (.A1(_11505_),
    .A2(_04273_),
    .A3(_04356_),
    .ZN(_04357_));
 AOI21_X4 _21348_ (.A(_04354_),
    .B1(_04355_),
    .B2(_04357_),
    .ZN(_04358_));
 BUF_X4 _21349_ (.A(_04358_),
    .Z(_04359_));
 CLKBUF_X3 _21350_ (.A(_04359_),
    .Z(_04360_));
 NOR3_X4 _21351_ (.A1(_04267_),
    .A2(_04354_),
    .A3(_04356_),
    .ZN(_04361_));
 BUF_X4 _21352_ (.A(_04361_),
    .Z(_04362_));
 CLKBUF_X3 _21353_ (.A(_04362_),
    .Z(_04363_));
 AOI22_X1 _21354_ (.A1(_16015_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_16018_),
    .ZN(_04364_));
 NOR2_X1 _21355_ (.A1(_04353_),
    .A2(_04364_),
    .ZN(_04365_));
 NOR2_X2 _21356_ (.A1(net301),
    .A2(_11505_),
    .ZN(_04366_));
 NOR3_X4 _21357_ (.A1(_04273_),
    .A2(_04354_),
    .A3(_04366_),
    .ZN(_04367_));
 BUF_X4 _21358_ (.A(_04367_),
    .Z(_04368_));
 BUF_X4 _21359_ (.A(_04368_),
    .Z(_04369_));
 CLKBUF_X3 _21360_ (.A(_04352_),
    .Z(_04370_));
 INV_X1 _21361_ (.A(_16014_),
    .ZN(_04371_));
 AOI221_X2 _21362_ (.A(_04365_),
    .B1(_04369_),
    .B2(\alu_adder_result_ex[22] ),
    .C1(_04370_),
    .C2(_04371_),
    .ZN(_04372_));
 AND3_X1 _21363_ (.A1(_15365_),
    .A2(_11482_),
    .A3(_11862_),
    .ZN(_04373_));
 AND3_X1 _21364_ (.A1(_11486_),
    .A2(_04264_),
    .A3(_11862_),
    .ZN(_04374_));
 MUX2_X2 _21365_ (.A(_04373_),
    .B(_04374_),
    .S(_11500_),
    .Z(_04375_));
 NAND2_X1 _21366_ (.A1(_04264_),
    .A2(_04273_),
    .ZN(_04376_));
 NOR2_X1 _21367_ (.A1(_04271_),
    .A2(_04269_),
    .ZN(_04377_));
 OAI22_X1 _21368_ (.A1(_04273_),
    .A2(_04304_),
    .B1(_04376_),
    .B2(_04377_),
    .ZN(_04378_));
 NAND2_X1 _21369_ (.A1(_04272_),
    .A2(_04268_),
    .ZN(_04379_));
 NOR2_X1 _21370_ (.A1(_04300_),
    .A2(_11512_),
    .ZN(_04380_));
 AOI221_X2 _21371_ (.A(_04375_),
    .B1(_04378_),
    .B2(_11862_),
    .C1(_04379_),
    .C2(_04380_),
    .ZN(_04381_));
 OAI21_X1 _21372_ (.A(_04268_),
    .B1(_04264_),
    .B2(_11476_),
    .ZN(_04382_));
 AOI22_X1 _21373_ (.A1(net301),
    .A2(_04376_),
    .B1(_04382_),
    .B2(_04267_),
    .ZN(_04383_));
 OR2_X1 _21374_ (.A1(_04265_),
    .A2(_04383_),
    .ZN(_04384_));
 NOR2_X1 _21375_ (.A1(net298),
    .A2(_04271_),
    .ZN(_04385_));
 OAI21_X1 _21376_ (.A(_04385_),
    .B1(_04366_),
    .B2(_04267_),
    .ZN(_04386_));
 NAND2_X2 _21377_ (.A1(_04348_),
    .A2(_04386_),
    .ZN(_04387_));
 NAND4_X2 _21378_ (.A1(_04381_),
    .A2(_04384_),
    .A3(_04387_),
    .A4(_04342_),
    .ZN(_04388_));
 NAND2_X1 _21379_ (.A1(_11406_),
    .A2(_04388_),
    .ZN(_04389_));
 BUF_X4 _21380_ (.A(_04389_),
    .Z(_04390_));
 BUF_X4 _21381_ (.A(_04390_),
    .Z(_04391_));
 OAI21_X2 _21382_ (.A(_04347_),
    .B1(_04372_),
    .B2(_04391_),
    .ZN(_04392_));
 BUF_X4 _21383_ (.A(_10744_),
    .Z(_04393_));
 NAND3_X1 _21384_ (.A1(_04316_),
    .A2(_04295_),
    .A3(_04343_),
    .ZN(_04394_));
 OAI21_X1 _21385_ (.A(_04305_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04395_));
 NAND3_X2 _21386_ (.A1(_15841_),
    .A2(_04394_),
    .A3(_04395_),
    .ZN(_04396_));
 CLKBUF_X3 _21387_ (.A(_10739_),
    .Z(_04397_));
 NAND4_X1 _21388_ (.A1(_04397_),
    .A2(_04316_),
    .A3(_04295_),
    .A4(_04314_),
    .ZN(_04398_));
 MUX2_X2 _21389_ (.A(_15838_),
    .B(_15492_),
    .S(_04302_),
    .Z(_04399_));
 OAI21_X1 _21390_ (.A(_04399_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04400_));
 AND3_X1 _21391_ (.A1(_04332_),
    .A2(_04398_),
    .A3(_04400_),
    .ZN(_04401_));
 OR2_X1 _21392_ (.A1(_10738_),
    .A2(_04321_),
    .ZN(_04402_));
 OAI21_X1 _21393_ (.A(_04402_),
    .B1(_04336_),
    .B2(_10739_),
    .ZN(_04403_));
 OR2_X1 _21394_ (.A1(_10739_),
    .A2(_04334_),
    .ZN(_04404_));
 OAI21_X1 _21395_ (.A(_04404_),
    .B1(_04327_),
    .B2(_15841_),
    .ZN(_04405_));
 NOR2_X4 _21396_ (.A1(_04318_),
    .A2(_04320_),
    .ZN(_04406_));
 MUX2_X1 _21397_ (.A(_04403_),
    .B(_04405_),
    .S(_04406_),
    .Z(_04407_));
 OR2_X1 _21398_ (.A1(_04297_),
    .A2(_04296_),
    .ZN(_04408_));
 BUF_X4 _21399_ (.A(_04408_),
    .Z(_04409_));
 BUF_X4 _21400_ (.A(_04409_),
    .Z(_04410_));
 AOI22_X4 _21401_ (.A1(_04396_),
    .A2(_04401_),
    .B1(_04407_),
    .B2(_04410_),
    .ZN(_04411_));
 NAND2_X4 _21402_ (.A1(_04279_),
    .A2(_04280_),
    .ZN(_04412_));
 NOR2_X1 _21403_ (.A1(_04412_),
    .A2(_04292_),
    .ZN(_04413_));
 NAND2_X1 _21404_ (.A1(_04411_),
    .A2(_04413_),
    .ZN(_04414_));
 MUX2_X1 _21405_ (.A(_15921_),
    .B(_16005_),
    .S(_04312_),
    .Z(_04415_));
 OR2_X1 _21406_ (.A1(_10738_),
    .A2(_04415_),
    .ZN(_04416_));
 OAI21_X1 _21407_ (.A(_04416_),
    .B1(_04325_),
    .B2(_10739_),
    .ZN(_04417_));
 MUX2_X1 _21408_ (.A(_15901_),
    .B(_16020_),
    .S(_04313_),
    .Z(_04418_));
 MUX2_X1 _21409_ (.A(_15893_),
    .B(_16033_),
    .S(_04313_),
    .Z(_04419_));
 MUX2_X1 _21410_ (.A(_04418_),
    .B(_04419_),
    .S(_10738_),
    .Z(_04420_));
 MUX2_X1 _21411_ (.A(_04417_),
    .B(_04420_),
    .S(_04330_),
    .Z(_04421_));
 MUX2_X1 _21412_ (.A(_15944_),
    .B(_15981_),
    .S(_04312_),
    .Z(_04422_));
 MUX2_X1 _21413_ (.A(_15952_),
    .B(_15976_),
    .S(_04312_),
    .Z(_04423_));
 MUX2_X1 _21414_ (.A(_04422_),
    .B(_04423_),
    .S(_10736_),
    .Z(_04424_));
 AND3_X1 _21415_ (.A1(_04315_),
    .A2(_04294_),
    .A3(_04424_),
    .ZN(_04425_));
 MUX2_X1 _21416_ (.A(_15928_),
    .B(_15997_),
    .S(_04312_),
    .Z(_04426_));
 MUX2_X1 _21417_ (.A(_15936_),
    .B(_15992_),
    .S(_04312_),
    .Z(_04427_));
 MUX2_X1 _21418_ (.A(_04426_),
    .B(_04427_),
    .S(_10739_),
    .Z(_04428_));
 BUF_X4 _21419_ (.A(_04330_),
    .Z(_04429_));
 AOI21_X1 _21420_ (.A(_04425_),
    .B1(_04428_),
    .B2(_04429_),
    .ZN(_04430_));
 BUF_X4 _21421_ (.A(_04409_),
    .Z(_04431_));
 MUX2_X1 _21422_ (.A(_04421_),
    .B(_04430_),
    .S(_04431_),
    .Z(_04432_));
 NOR2_X4 _21423_ (.A1(net278),
    .A2(_04310_),
    .ZN(_04433_));
 CLKBUF_X3 _21424_ (.A(_04433_),
    .Z(_04434_));
 XNOR2_X1 _21425_ (.A(_10739_),
    .B(_04434_),
    .ZN(_04435_));
 MUX2_X1 _21426_ (.A(_15961_),
    .B(_15964_),
    .S(_04435_),
    .Z(_04436_));
 MUX2_X1 _21427_ (.A(_15952_),
    .B(_15976_),
    .S(_04433_),
    .Z(_04437_));
 MUX2_X1 _21428_ (.A(_15944_),
    .B(_15981_),
    .S(_04433_),
    .Z(_04438_));
 MUX2_X1 _21429_ (.A(_04437_),
    .B(_04438_),
    .S(_10739_),
    .Z(_04439_));
 INV_X1 _21430_ (.A(_04439_),
    .ZN(_04440_));
 MUX2_X1 _21431_ (.A(_04436_),
    .B(_04440_),
    .S(_04406_),
    .Z(_04441_));
 MUX2_X1 _21432_ (.A(_15921_),
    .B(_16005_),
    .S(_04433_),
    .Z(_04442_));
 OR2_X1 _21433_ (.A1(_04397_),
    .A2(_04442_),
    .ZN(_04443_));
 MUX2_X1 _21434_ (.A(_15913_),
    .B(_16013_),
    .S(_04434_),
    .Z(_04444_));
 OAI21_X1 _21435_ (.A(_04443_),
    .B1(_04444_),
    .B2(_15841_),
    .ZN(_04445_));
 MUX2_X1 _21436_ (.A(_15936_),
    .B(_15992_),
    .S(_04433_),
    .Z(_04446_));
 MUX2_X1 _21437_ (.A(_15928_),
    .B(_15997_),
    .S(_04433_),
    .Z(_04447_));
 MUX2_X1 _21438_ (.A(_04446_),
    .B(_04447_),
    .S(_10739_),
    .Z(_04448_));
 INV_X1 _21439_ (.A(_04448_),
    .ZN(_04449_));
 MUX2_X1 _21440_ (.A(_04445_),
    .B(_04449_),
    .S(_04429_),
    .Z(_04450_));
 MUX2_X1 _21441_ (.A(_04441_),
    .B(_04450_),
    .S(_04431_),
    .Z(_04451_));
 NAND2_X4 _21442_ (.A1(_04284_),
    .A2(_04290_),
    .ZN(_04452_));
 CLKBUF_X3 _21443_ (.A(_04452_),
    .Z(_04453_));
 MUX2_X1 _21444_ (.A(_04432_),
    .B(_04451_),
    .S(_04453_),
    .Z(_04454_));
 OAI21_X1 _21445_ (.A(_04414_),
    .B1(_04454_),
    .B2(_04308_),
    .ZN(_04455_));
 AND3_X2 _21446_ (.A1(_04271_),
    .A2(_04300_),
    .A3(_04301_),
    .ZN(_04456_));
 CLKBUF_X3 _21447_ (.A(_04456_),
    .Z(_04457_));
 NOR2_X2 _21448_ (.A1(_04452_),
    .A2(_04306_),
    .ZN(_04458_));
 NAND2_X1 _21449_ (.A1(_04281_),
    .A2(_04458_),
    .ZN(_04459_));
 NAND2_X1 _21450_ (.A1(_04457_),
    .A2(_04459_),
    .ZN(_04460_));
 XNOR2_X2 _21451_ (.A(_14125_),
    .B(_15619_),
    .ZN(_04461_));
 OR3_X1 _21452_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A2(_11430_),
    .A3(_11433_),
    .ZN(_04462_));
 CLKBUF_X3 _21453_ (.A(_04462_),
    .Z(_04463_));
 NOR2_X1 _21454_ (.A1(_04461_),
    .A2(_04463_),
    .ZN(_04464_));
 INV_X1 _21455_ (.A(_15757_),
    .ZN(_04465_));
 NOR2_X1 _21456_ (.A1(_15745_),
    .A2(_15744_),
    .ZN(_04466_));
 INV_X1 _21457_ (.A(_04466_),
    .ZN(_04467_));
 AOI21_X1 _21458_ (.A(_15750_),
    .B1(_04467_),
    .B2(_15751_),
    .ZN(_04468_));
 NOR2_X1 _21459_ (.A1(_04465_),
    .A2(_04468_),
    .ZN(_04469_));
 OAI21_X1 _21460_ (.A(_15763_),
    .B1(_15756_),
    .B2(_04469_),
    .ZN(_04470_));
 NOR4_X2 _21461_ (.A1(_15738_),
    .A2(_15744_),
    .A3(_15750_),
    .A4(_15756_),
    .ZN(_04471_));
 BUF_X4 _21462_ (.A(_15739_),
    .Z(_04472_));
 AND3_X2 _21463_ (.A1(_04472_),
    .A2(_15730_),
    .A3(_15726_),
    .ZN(_04473_));
 OR3_X4 _21464_ (.A1(_15716_),
    .A2(_15706_),
    .A3(_15699_),
    .ZN(_04474_));
 AOI21_X2 clone77 (.A(_03674_),
    .B1(_10470_),
    .B2(_10474_),
    .ZN(net348));
 OR3_X4 _21466_ (.A1(_15657_),
    .A2(_15671_),
    .A3(_15685_),
    .ZN(_04476_));
 INV_X1 _21467_ (.A(_15630_),
    .ZN(_04477_));
 AOI21_X1 _21468_ (.A(_15618_),
    .B1(_15619_),
    .B2(_14125_),
    .ZN(_04478_));
 INV_X1 _21469_ (.A(_15631_),
    .ZN(_04479_));
 OAI21_X2 _21470_ (.A(_04477_),
    .B1(_04478_),
    .B2(_04479_),
    .ZN(_04480_));
 BUF_X2 _21471_ (.A(_15644_),
    .Z(_04481_));
 AOI211_X2 _21472_ (.A(_15643_),
    .B(_04476_),
    .C1(_04480_),
    .C2(_04481_),
    .ZN(_04482_));
 BUF_X4 clone50 (.A(net322),
    .Z(net321));
 INV_X1 _21474_ (.A(_15686_),
    .ZN(_04484_));
 INV_X1 _21475_ (.A(_15671_),
    .ZN(_04485_));
 BUF_X2 _21476_ (.A(_15672_),
    .Z(_04486_));
 OAI21_X1 _21477_ (.A(_04486_),
    .B1(_15657_),
    .B2(_15658_),
    .ZN(_04487_));
 AOI21_X2 _21478_ (.A(_04484_),
    .B1(_04485_),
    .B2(_04487_),
    .ZN(_04488_));
 OAI21_X2 _21479_ (.A(_15700_),
    .B1(_15685_),
    .B2(_04488_),
    .ZN(_04489_));
 NOR2_X2 _21480_ (.A1(_04482_),
    .A2(_04489_),
    .ZN(_04490_));
 BUF_X2 _21481_ (.A(_15707_),
    .Z(_04491_));
 OAI21_X2 _21482_ (.A(_15717_),
    .B1(_15706_),
    .B2(_04491_),
    .ZN(_04492_));
 INV_X1 _21483_ (.A(_04492_),
    .ZN(_04493_));
 OAI221_X2 _21484_ (.A(_04473_),
    .B1(_04474_),
    .B2(_04490_),
    .C1(_15716_),
    .C2(_04493_),
    .ZN(_04494_));
 AOI21_X4 _21485_ (.A(_15729_),
    .B1(net318),
    .B2(_15725_),
    .ZN(_04495_));
 INV_X1 _21486_ (.A(_04495_),
    .ZN(_04496_));
 NAND2_X1 _21487_ (.A1(_04472_),
    .A2(_04496_),
    .ZN(_04497_));
 AND2_X4 _21488_ (.A1(_04494_),
    .A2(_04497_),
    .ZN(_04498_));
 AOI21_X4 _21489_ (.A(_04470_),
    .B1(_04498_),
    .B2(_04471_),
    .ZN(_04499_));
 NOR2_X1 _21490_ (.A1(_15762_),
    .A2(_04499_),
    .ZN(_04500_));
 XNOR2_X1 _21491_ (.A(_15769_),
    .B(_04500_),
    .ZN(_04501_));
 CLKBUF_X3 _21492_ (.A(_04463_),
    .Z(_04502_));
 AOI21_X2 _21493_ (.A(_04464_),
    .B1(_04501_),
    .B2(_04502_),
    .ZN(_04503_));
 MUX2_X2 _21494_ (.A(_03813_),
    .B(_04503_),
    .S(_12102_),
    .Z(_04504_));
 OAI221_X2 _21495_ (.A(_04393_),
    .B1(_04455_),
    .B2(_04460_),
    .C1(_04504_),
    .C2(_11408_),
    .ZN(_04505_));
 NAND3_X2 _21496_ (.A1(_10921_),
    .A2(_15888_),
    .A3(_15892_),
    .ZN(_04506_));
 OAI21_X2 _21497_ (.A(_11116_),
    .B1(_11063_),
    .B2(_11061_),
    .ZN(_04507_));
 OR4_X1 _21498_ (.A1(_15920_),
    .A2(_04238_),
    .A3(_04506_),
    .A4(_04507_),
    .ZN(_04508_));
 BUF_X4 _21499_ (.A(_04508_),
    .Z(_04509_));
 AOI211_X2 _21500_ (.A(_03504_),
    .B(_04509_),
    .C1(_03540_),
    .C2(_10921_),
    .ZN(_04510_));
 BUF_X4 _21501_ (.A(net16),
    .Z(_04511_));
 NAND4_X4 _21502_ (.A1(_15929_),
    .A2(_03491_),
    .A3(_04248_),
    .A4(_03587_),
    .ZN(_04512_));
 NOR2_X1 _21503_ (.A1(_10920_),
    .A2(_03537_),
    .ZN(_04513_));
 NOR3_X4 _21504_ (.A1(_03575_),
    .A2(_04512_),
    .A3(_04513_),
    .ZN(_04514_));
 BUF_X4 _21505_ (.A(_04514_),
    .Z(_04515_));
 AOI22_X1 _21506_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_04511_),
    .B1(_04515_),
    .B2(\cs_registers_i.mie_q[6] ),
    .ZN(_04516_));
 NOR2_X4 _21507_ (.A1(_03575_),
    .A2(_04244_),
    .ZN(_04517_));
 BUF_X4 _21508_ (.A(_04517_),
    .Z(_04518_));
 AOI21_X2 _21509_ (.A(_04244_),
    .B1(_03577_),
    .B2(_03576_),
    .ZN(_04519_));
 BUF_X4 _21510_ (.A(_04519_),
    .Z(_04520_));
 BUF_X4 _21511_ (.A(_04520_),
    .Z(_04521_));
 AOI211_X2 _21512_ (.A(_03500_),
    .B(_04244_),
    .C1(_03518_),
    .C2(_03540_),
    .ZN(_04522_));
 BUF_X4 _21513_ (.A(_04522_),
    .Z(_04523_));
 BUF_X4 _21514_ (.A(_04523_),
    .Z(_04524_));
 AOI222_X2 _21515_ (.A1(net147),
    .A2(_04518_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[22] ),
    .C1(\cs_registers_i.mscratch_q[22] ),
    .C2(_04524_),
    .ZN(_04525_));
 AND3_X4 _21516_ (.A1(_03514_),
    .A2(_04255_),
    .A3(_03595_),
    .ZN(_04526_));
 BUF_X4 _21517_ (.A(_04526_),
    .Z(_04527_));
 BUF_X4 _21518_ (.A(_04527_),
    .Z(_04528_));
 AOI21_X4 _21519_ (.A(_04509_),
    .B1(_03576_),
    .B2(_03577_),
    .ZN(_04529_));
 BUF_X4 _21520_ (.A(_04529_),
    .Z(_04530_));
 AOI22_X1 _21521_ (.A1(net85),
    .A2(_04528_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[22] ),
    .ZN(_04531_));
 OR3_X1 _21522_ (.A1(_03580_),
    .A2(_03581_),
    .A3(_04512_),
    .ZN(_04532_));
 CLKBUF_X3 _21523_ (.A(_04532_),
    .Z(_04533_));
 BUF_X4 _21524_ (.A(_04533_),
    .Z(_04534_));
 NOR3_X4 _21525_ (.A1(_03502_),
    .A2(_10919_),
    .A3(_15876_),
    .ZN(_04535_));
 NAND4_X4 _21526_ (.A1(_15873_),
    .A2(_03594_),
    .A3(_04249_),
    .A4(_04535_),
    .ZN(_04536_));
 BUF_X4 _21527_ (.A(_04536_),
    .Z(_04537_));
 NOR4_X4 _21528_ (.A1(_15920_),
    .A2(_04238_),
    .A3(_04506_),
    .A4(_04507_),
    .ZN(_04538_));
 OAI211_X4 _21529_ (.A(_03501_),
    .B(_04538_),
    .C1(_03530_),
    .C2(_10920_),
    .ZN(_04539_));
 INV_X1 _21530_ (.A(\cs_registers_i.csr_depc_o[22] ),
    .ZN(_04540_));
 OAI221_X2 _21531_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01179_),
    .C1(_04539_),
    .C2(_04540_),
    .ZN(_04541_));
 AOI211_X2 _21532_ (.A(_03502_),
    .B(_04244_),
    .C1(_03540_),
    .C2(_10922_),
    .ZN(_04542_));
 BUF_X4 _21533_ (.A(_04542_),
    .Z(_04543_));
 BUF_X4 _21534_ (.A(_04543_),
    .Z(_04544_));
 AOI21_X2 _21535_ (.A(_04541_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[22] ),
    .ZN(_04545_));
 AND4_X1 _21536_ (.A1(_04516_),
    .A2(_04525_),
    .A3(_04531_),
    .A4(_04545_),
    .ZN(_04546_));
 BUF_X2 _21537_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .Z(_04547_));
 OR4_X2 _21538_ (.A1(_15508_),
    .A2(_03501_),
    .A3(_03506_),
    .A4(_03503_),
    .ZN(_04548_));
 AOI21_X4 _21539_ (.A(_04548_),
    .B1(_03574_),
    .B2(_03540_),
    .ZN(_04549_));
 BUF_X4 _21540_ (.A(_04549_),
    .Z(_04550_));
 BUF_X4 _21541_ (.A(_04550_),
    .Z(_04551_));
 AOI21_X4 _21542_ (.A(_03504_),
    .B1(_10922_),
    .B2(_03580_),
    .ZN(_04552_));
 BUF_X4 _21543_ (.A(_04552_),
    .Z(_04553_));
 BUF_X4 _21544_ (.A(_04553_),
    .Z(_04554_));
 AOI22_X2 _21545_ (.A1(_04547_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][54] ),
    .ZN(_04555_));
 OR2_X1 _21546_ (.A1(_03551_),
    .A2(_04236_),
    .ZN(_04556_));
 BUF_X4 _21547_ (.A(_04556_),
    .Z(_04557_));
 BUF_X4 _21548_ (.A(_04557_),
    .Z(_04558_));
 CLKBUF_X3 _21549_ (.A(_04235_),
    .Z(_04559_));
 BUF_X4 _21550_ (.A(_04559_),
    .Z(_04560_));
 AOI22_X2 _21551_ (.A1(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][22] ),
    .ZN(_04561_));
 OAI221_X2 _21552_ (.A(_04546_),
    .B1(_04555_),
    .B2(_04558_),
    .C1(_04560_),
    .C2(_04561_),
    .ZN(_04562_));
 BUF_X4 _21553_ (.A(_04393_),
    .Z(_04563_));
 OAI221_X2 _21554_ (.A(_04263_),
    .B1(_04505_),
    .B2(_04392_),
    .C1(_04562_),
    .C2(_04563_),
    .ZN(_04564_));
 BUF_X4 _21555_ (.A(\load_store_unit_i.data_type_q[1] ),
    .Z(_04565_));
 CLKBUF_X2 _21556_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_04566_));
 MUX2_X1 _21557_ (.A(net66),
    .B(net44),
    .S(_04566_),
    .Z(_04567_));
 BUF_X1 _21558_ (.A(data_rdata_i[23]),
    .Z(_04568_));
 MUX2_X1 _21559_ (.A(_04568_),
    .B(net61),
    .S(_04566_),
    .Z(_04569_));
 BUF_X4 _21560_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_04570_));
 MUX2_X1 _21561_ (.A(_04567_),
    .B(_04569_),
    .S(_04570_),
    .Z(_04571_));
 NAND3_X4 _21562_ (.A1(_04565_),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_04571_),
    .ZN(_04572_));
 BUF_X2 _21563_ (.A(\load_store_unit_i.data_type_q[2] ),
    .Z(_04573_));
 BUF_X4 _21564_ (.A(_04573_),
    .Z(_04574_));
 MUX2_X1 _21565_ (.A(net61),
    .B(net66),
    .S(_04566_),
    .Z(_04575_));
 MUX2_X1 _21566_ (.A(net44),
    .B(_04568_),
    .S(_04566_),
    .Z(_04576_));
 INV_X2 _21567_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .ZN(_04577_));
 MUX2_X1 _21568_ (.A(_04575_),
    .B(_04576_),
    .S(_04577_),
    .Z(_04578_));
 NAND3_X2 _21569_ (.A1(_04574_),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_04578_),
    .ZN(_04579_));
 NAND2_X4 _21570_ (.A1(_04572_),
    .A2(_04579_),
    .ZN(_04580_));
 NOR2_X4 _21571_ (.A1(_04573_),
    .A2(_04565_),
    .ZN(_04581_));
 BUF_X4 _21572_ (.A(_04581_),
    .Z(_04582_));
 BUF_X4 _21573_ (.A(_04582_),
    .Z(_04583_));
 BUF_X4 _21574_ (.A(_04566_),
    .Z(_04584_));
 CLKBUF_X3 _21575_ (.A(_04584_),
    .Z(_04585_));
 CLKBUF_X3 _21576_ (.A(_04585_),
    .Z(_04586_));
 NOR2_X1 _21577_ (.A1(_04586_),
    .A2(net65),
    .ZN(_04587_));
 INV_X1 _21578_ (.A(_04566_),
    .ZN(_04588_));
 CLKBUF_X3 _21579_ (.A(_04588_),
    .Z(_04589_));
 NOR2_X1 _21580_ (.A1(_04589_),
    .A2(net43),
    .ZN(_04590_));
 OR3_X1 _21581_ (.A1(_04577_),
    .A2(_04587_),
    .A3(_04590_),
    .ZN(_04591_));
 AND2_X1 _21582_ (.A1(_04588_),
    .A2(net52),
    .ZN(_04592_));
 CLKBUF_X3 _21583_ (.A(_04584_),
    .Z(_04593_));
 BUF_X4 _21584_ (.A(_04593_),
    .Z(_04594_));
 AOI21_X1 _21585_ (.A(_04592_),
    .B1(\load_store_unit_i.rdata_q[30] ),
    .B2(_04594_),
    .ZN(_04595_));
 CLKBUF_X3 _21586_ (.A(_04570_),
    .Z(_04596_));
 BUF_X4 _21587_ (.A(_04596_),
    .Z(_04597_));
 OAI21_X1 _21588_ (.A(_04591_),
    .B1(_04595_),
    .B2(_04597_),
    .ZN(_04598_));
 AOI21_X2 _21589_ (.A(_04580_),
    .B1(_04583_),
    .B2(_04598_),
    .ZN(_04599_));
 BUF_X8 _21590_ (.A(_04263_),
    .Z(_04600_));
 OAI21_X4 _21591_ (.A(_04564_),
    .B1(_04599_),
    .B2(_04600_),
    .ZN(_04601_));
 BUF_X2 _21592_ (.A(_04601_),
    .Z(_04602_));
 BUF_X4 _21593_ (.A(_00039_),
    .Z(_04603_));
 NOR3_X4 _21594_ (.A1(_10394_),
    .A2(_11315_),
    .A3(_04603_),
    .ZN(_04604_));
 NAND4_X4 _21595_ (.A1(_03453_),
    .A2(_01160_),
    .A3(_03455_),
    .A4(_03457_),
    .ZN(_04605_));
 NOR4_X2 _21596_ (.A1(_03518_),
    .A2(_11428_),
    .A3(_04229_),
    .A4(_04231_),
    .ZN(_04606_));
 NOR4_X4 _21597_ (.A1(_11428_),
    .A2(_03508_),
    .A3(_04229_),
    .A4(_04231_),
    .ZN(_04607_));
 OAI21_X1 _21598_ (.A(_03532_),
    .B1(_03536_),
    .B2(_03551_),
    .ZN(_04608_));
 OR2_X1 _21599_ (.A1(_03603_),
    .A2(_04608_),
    .ZN(_04609_));
 AOI21_X4 _21600_ (.A(_04606_),
    .B1(_04607_),
    .B2(_04609_),
    .ZN(_04610_));
 BUF_X4 _21601_ (.A(_04610_),
    .Z(_04611_));
 AOI211_X2 _21602_ (.A(_10900_),
    .B(_10901_),
    .C1(_04605_),
    .C2(_04611_),
    .ZN(_04612_));
 BUF_X8 _21603_ (.A(_04612_),
    .Z(_04613_));
 NAND2_X4 _21604_ (.A1(_04604_),
    .A2(_04613_),
    .ZN(_04614_));
 BUF_X4 _21605_ (.A(_04614_),
    .Z(_04615_));
 MUX2_X1 _21606_ (.A(_04602_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .S(_04615_),
    .Z(_01185_));
 INV_X1 _21607_ (.A(_04580_),
    .ZN(_04616_));
 NAND2_X4 _21608_ (.A1(_04611_),
    .A2(_04616_),
    .ZN(_04617_));
 MUX2_X1 _21609_ (.A(_04568_),
    .B(\load_store_unit_i.rdata_q[31] ),
    .S(_04593_),
    .Z(_04618_));
 CLKBUF_X3 _21610_ (.A(_04577_),
    .Z(_04619_));
 MUX2_X1 _21611_ (.A(_04567_),
    .B(_04618_),
    .S(_04619_),
    .Z(_04620_));
 AOI21_X2 _21612_ (.A(_04617_),
    .B1(_04620_),
    .B2(_04583_),
    .ZN(_04621_));
 BUF_X4 _21613_ (.A(_10493_),
    .Z(_04622_));
 NOR3_X2 _21614_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A2(_11430_),
    .A3(_11433_),
    .ZN(_04623_));
 CLKBUF_X3 _21615_ (.A(_04623_),
    .Z(_04624_));
 CLKBUF_X3 _21616_ (.A(_04624_),
    .Z(_04625_));
 CLKBUF_X3 _21617_ (.A(_04625_),
    .Z(_04626_));
 INV_X1 _21618_ (.A(_15618_),
    .ZN(_04627_));
 AOI21_X1 _21619_ (.A(_15599_),
    .B1(_15600_),
    .B2(_14124_),
    .ZN(_04628_));
 INV_X1 _21620_ (.A(_15619_),
    .ZN(_04629_));
 OAI21_X2 _21621_ (.A(_04627_),
    .B1(_04628_),
    .B2(_04629_),
    .ZN(_04630_));
 XNOR2_X2 _21622_ (.A(_04479_),
    .B(_04630_),
    .ZN(_04631_));
 AOI21_X1 _21623_ (.A(_04622_),
    .B1(_04626_),
    .B2(_04631_),
    .ZN(_04632_));
 INV_X1 _21624_ (.A(_15763_),
    .ZN(_04633_));
 INV_X1 _21625_ (.A(_15756_),
    .ZN(_04634_));
 INV_X1 _21626_ (.A(_15750_),
    .ZN(_04635_));
 NOR2_X1 _21627_ (.A1(_15738_),
    .A2(_15744_),
    .ZN(_04636_));
 NAND2_X1 _21628_ (.A1(_04635_),
    .A2(_04636_),
    .ZN(_04637_));
 NAND2_X2 _21629_ (.A1(_15726_),
    .A2(_15730_),
    .ZN(_04638_));
 INV_X1 _21630_ (.A(_15716_),
    .ZN(_04639_));
 AOI21_X4 _21631_ (.A(_04638_),
    .B1(_04492_),
    .B2(_04639_),
    .ZN(_04640_));
 AND2_X1 _21632_ (.A1(_15700_),
    .A2(_15685_),
    .ZN(_04641_));
 OR2_X4 _21633_ (.A1(_04474_),
    .A2(_04641_),
    .ZN(_04642_));
 NAND3_X4 _21634_ (.A1(_04472_),
    .A2(_04640_),
    .A3(_04642_),
    .ZN(_04643_));
 NAND2_X4 _21635_ (.A1(_04497_),
    .A2(_04643_),
    .ZN(_04644_));
 AND3_X4 _21636_ (.A1(_15700_),
    .A2(_04472_),
    .A3(_04640_),
    .ZN(_04645_));
 INV_X2 _21637_ (.A(_04486_),
    .ZN(_04646_));
 AOI21_X1 _21638_ (.A(_15657_),
    .B1(_15643_),
    .B2(_15658_),
    .ZN(_04647_));
 NOR2_X1 _21639_ (.A1(_04646_),
    .A2(_04647_),
    .ZN(_04648_));
 OAI21_X2 _21640_ (.A(_15686_),
    .B1(_15671_),
    .B2(_04648_),
    .ZN(_04649_));
 AOI21_X4 _21641_ (.A(_15630_),
    .B1(_04630_),
    .B2(_15631_),
    .ZN(_04650_));
 NAND4_X1 _21642_ (.A1(_04481_),
    .A2(_15658_),
    .A3(_04486_),
    .A4(_15686_),
    .ZN(_04651_));
 OAI21_X2 _21643_ (.A(_04649_),
    .B1(_04650_),
    .B2(_04651_),
    .ZN(_04652_));
 AOI211_X2 _21644_ (.A(_04637_),
    .B(_04644_),
    .C1(_04645_),
    .C2(_04652_),
    .ZN(_04653_));
 OR3_X4 _21645_ (.A1(_04653_),
    .A2(_04468_),
    .A3(_04465_),
    .ZN(_04654_));
 AOI21_X4 _21646_ (.A(_04633_),
    .B1(_04654_),
    .B2(_04634_),
    .ZN(_04655_));
 OR2_X1 _21647_ (.A1(_15762_),
    .A2(_04655_),
    .ZN(_04656_));
 AOI21_X1 _21648_ (.A(_15768_),
    .B1(_04656_),
    .B2(_15769_),
    .ZN(_04657_));
 XOR2_X1 _21649_ (.A(_15775_),
    .B(_04657_),
    .Z(_04658_));
 OAI21_X1 _21650_ (.A(_04632_),
    .B1(_04658_),
    .B2(_04626_),
    .ZN(_04659_));
 AOI21_X1 _21651_ (.A(_11408_),
    .B1(_03815_),
    .B2(net300),
    .ZN(_04660_));
 AND2_X2 _21652_ (.A1(_04659_),
    .A2(_04660_),
    .ZN(_04661_));
 BUF_X8 _21653_ (.A(_03493_),
    .Z(_04662_));
 AOI22_X1 _21654_ (.A1(_16023_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_16022_),
    .ZN(_04663_));
 NAND2_X4 _21655_ (.A1(_04348_),
    .A2(_04349_),
    .ZN(_04664_));
 CLKBUF_X3 _21656_ (.A(_04664_),
    .Z(_04665_));
 MUX2_X1 _21657_ (.A(_16026_),
    .B(_04663_),
    .S(_04665_),
    .Z(_04666_));
 NAND2_X1 _21658_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_04369_),
    .ZN(_04667_));
 AOI21_X1 _21659_ (.A(_04390_),
    .B1(_04666_),
    .B2(_04667_),
    .ZN(_04668_));
 NOR2_X1 _21660_ (.A1(_04662_),
    .A2(_04668_),
    .ZN(_04669_));
 NAND2_X2 _21661_ (.A1(_04412_),
    .A2(_04292_),
    .ZN(_04670_));
 INV_X1 _21662_ (.A(_11497_),
    .ZN(_04671_));
 OR4_X1 _21663_ (.A1(_04671_),
    .A2(_04304_),
    .A3(_04265_),
    .A4(_04399_),
    .ZN(_04672_));
 NOR2_X2 _21664_ (.A1(_04409_),
    .A2(_04672_),
    .ZN(_04673_));
 NAND2_X2 _21665_ (.A1(_04303_),
    .A2(_04305_),
    .ZN(_04674_));
 NAND3_X1 _21666_ (.A1(_04397_),
    .A2(_04316_),
    .A3(_04295_),
    .ZN(_04675_));
 OAI21_X2 _21667_ (.A(_04674_),
    .B1(_04675_),
    .B2(_04399_),
    .ZN(_04676_));
 AOI21_X2 _21668_ (.A(_04673_),
    .B1(_04676_),
    .B2(_04431_),
    .ZN(_04677_));
 NOR2_X2 _21669_ (.A1(_04670_),
    .A2(_04677_),
    .ZN(_04678_));
 OR2_X1 _21670_ (.A1(_04322_),
    .A2(_04317_),
    .ZN(_04679_));
 MUX2_X1 _21671_ (.A(_15865_),
    .B(_16060_),
    .S(_04302_),
    .Z(_04680_));
 MUX2_X1 _21672_ (.A(_04680_),
    .B(_04343_),
    .S(_04330_),
    .Z(_04681_));
 MUX2_X1 _21673_ (.A(_04679_),
    .B(_04681_),
    .S(_15841_),
    .Z(_04682_));
 MUX2_X1 _21674_ (.A(_04420_),
    .B(_04405_),
    .S(_04429_),
    .Z(_04683_));
 MUX2_X2 _21675_ (.A(_04682_),
    .B(_04683_),
    .S(_04410_),
    .Z(_04684_));
 AOI22_X4 _21676_ (.A1(_04279_),
    .A2(_04280_),
    .B1(_04284_),
    .B2(_04290_),
    .ZN(_04685_));
 AOI221_X2 _21677_ (.A(_04678_),
    .B1(_04684_),
    .B2(_04685_),
    .C1(_04282_),
    .C2(_04307_),
    .ZN(_04686_));
 OR4_X4 _21678_ (.A1(_04264_),
    .A2(_04265_),
    .A3(_04270_),
    .A4(_04274_),
    .ZN(_04687_));
 BUF_X4 _21679_ (.A(_04687_),
    .Z(_04688_));
 MUX2_X1 _21680_ (.A(_15852_),
    .B(_16068_),
    .S(_04313_),
    .Z(_04689_));
 MUX2_X1 _21681_ (.A(_04689_),
    .B(_04680_),
    .S(_10739_),
    .Z(_04690_));
 MUX2_X2 _21682_ (.A(_04344_),
    .B(_04690_),
    .S(_04406_),
    .Z(_04691_));
 NAND2_X2 _21683_ (.A1(_04406_),
    .A2(_04329_),
    .ZN(_04692_));
 MUX2_X1 _21684_ (.A(_04321_),
    .B(_04334_),
    .S(_10739_),
    .Z(_04693_));
 AOI21_X2 _21685_ (.A(_04332_),
    .B1(_04429_),
    .B2(_04693_),
    .ZN(_04694_));
 AOI22_X4 _21686_ (.A1(_04333_),
    .A2(_04691_),
    .B1(_04692_),
    .B2(_04694_),
    .ZN(_04695_));
 AOI211_X2 _21687_ (.A(_04412_),
    .B(_04458_),
    .C1(_04695_),
    .C2(_04453_),
    .ZN(_04696_));
 MUX2_X1 _21688_ (.A(_04415_),
    .B(_04426_),
    .S(_10739_),
    .Z(_04697_));
 AND3_X1 _21689_ (.A1(_04316_),
    .A2(_04295_),
    .A3(_04697_),
    .ZN(_04698_));
 AOI21_X2 _21690_ (.A(_04698_),
    .B1(_04326_),
    .B2(_04429_),
    .ZN(_04699_));
 MUX2_X1 _21691_ (.A(_15957_),
    .B(_15968_),
    .S(_04313_),
    .Z(_04700_));
 MUX2_X1 _21692_ (.A(_04423_),
    .B(_04700_),
    .S(_04397_),
    .Z(_04701_));
 NAND3_X1 _21693_ (.A1(_04316_),
    .A2(_04295_),
    .A3(_04701_),
    .ZN(_04702_));
 MUX2_X1 _21694_ (.A(_04422_),
    .B(_04427_),
    .S(_10738_),
    .Z(_04703_));
 OAI21_X1 _21695_ (.A(_04703_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04704_));
 AND2_X1 _21696_ (.A1(_04702_),
    .A2(_04704_),
    .ZN(_04705_));
 MUX2_X1 _21697_ (.A(_04699_),
    .B(_04705_),
    .S(_04431_),
    .Z(_04706_));
 CLKBUF_X3 _21698_ (.A(_04410_),
    .Z(_04707_));
 MUX2_X1 _21699_ (.A(_04438_),
    .B(_04446_),
    .S(_10739_),
    .Z(_04708_));
 MUX2_X1 _21700_ (.A(_15957_),
    .B(_15968_),
    .S(_04433_),
    .Z(_04709_));
 MUX2_X1 _21701_ (.A(_04437_),
    .B(_04709_),
    .S(_10738_),
    .Z(_04710_));
 MUX2_X1 _21702_ (.A(_04708_),
    .B(_04710_),
    .S(_04429_),
    .Z(_04711_));
 CLKBUF_X3 _21703_ (.A(_04406_),
    .Z(_04712_));
 MUX2_X1 _21704_ (.A(_15905_),
    .B(_16024_),
    .S(_04434_),
    .Z(_04713_));
 MUX2_X1 _21705_ (.A(_04444_),
    .B(_04713_),
    .S(_04397_),
    .Z(_04714_));
 AND2_X1 _21706_ (.A1(_04712_),
    .A2(_04714_),
    .ZN(_04715_));
 MUX2_X1 _21707_ (.A(_04442_),
    .B(_04447_),
    .S(_10738_),
    .Z(_04716_));
 OAI21_X1 _21708_ (.A(_04716_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04717_));
 NAND2_X1 _21709_ (.A1(_04431_),
    .A2(_04717_),
    .ZN(_04718_));
 OAI22_X1 _21710_ (.A1(_04707_),
    .A2(_04711_),
    .B1(_04715_),
    .B2(_04718_),
    .ZN(_04719_));
 CLKBUF_X3 _21711_ (.A(_04453_),
    .Z(_04720_));
 MUX2_X1 _21712_ (.A(_04706_),
    .B(_04719_),
    .S(_04720_),
    .Z(_04721_));
 CLKBUF_X3 _21713_ (.A(_04412_),
    .Z(_04722_));
 BUF_X4 _21714_ (.A(_04722_),
    .Z(_04723_));
 AOI21_X2 _21715_ (.A(_04696_),
    .B1(_04721_),
    .B2(_04723_),
    .ZN(_04724_));
 BUF_X4 _21716_ (.A(_04302_),
    .Z(_04725_));
 OAI221_X2 _21717_ (.A(_04669_),
    .B1(_04686_),
    .B2(_04688_),
    .C1(_04724_),
    .C2(_04725_),
    .ZN(_04726_));
 AND3_X1 _21718_ (.A1(_03501_),
    .A2(_15873_),
    .A3(_03570_),
    .ZN(_04727_));
 NAND3_X2 _21719_ (.A1(_03594_),
    .A2(_03588_),
    .A3(_04727_),
    .ZN(_04728_));
 NOR2_X1 _21720_ (.A1(_01180_),
    .A2(_04728_),
    .ZN(_04729_));
 OAI21_X2 _21721_ (.A(_03503_),
    .B1(_03530_),
    .B2(_03499_),
    .ZN(_04730_));
 NOR2_X4 _21722_ (.A1(_03498_),
    .A2(_04730_),
    .ZN(_04731_));
 OAI21_X2 _21723_ (.A(_03588_),
    .B1(_03537_),
    .B2(_03499_),
    .ZN(_04732_));
 NOR2_X4 _21724_ (.A1(_03575_),
    .A2(_04732_),
    .ZN(_04733_));
 AOI221_X2 _21725_ (.A(_04729_),
    .B1(_04731_),
    .B2(\cs_registers_i.dscratch0_q[23] ),
    .C1(\cs_registers_i.mie_q[7] ),
    .C2(_04733_),
    .ZN(_04734_));
 OAI21_X4 _21726_ (.A(_03501_),
    .B1(_10920_),
    .B2(_03530_),
    .ZN(_04735_));
 NOR2_X4 _21727_ (.A1(_03498_),
    .A2(_04735_),
    .ZN(_04736_));
 NAND2_X4 _21728_ (.A1(_03553_),
    .A2(_03572_),
    .ZN(_04737_));
 NOR2_X2 _21729_ (.A1(_11072_),
    .A2(_04737_),
    .ZN(_04738_));
 AOI22_X2 _21730_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_04736_),
    .B1(_04738_),
    .B2(\cs_registers_i.mscratch_q[23] ),
    .ZN(_04739_));
 NOR2_X1 _21731_ (.A1(_03580_),
    .A2(_03581_),
    .ZN(_04740_));
 AND2_X2 _21732_ (.A1(_04740_),
    .A2(_03588_),
    .ZN(_04741_));
 NOR2_X2 _21733_ (.A1(_03575_),
    .A2(_04737_),
    .ZN(_04742_));
 AND4_X2 _21734_ (.A1(_03564_),
    .A2(_03594_),
    .A3(_03595_),
    .A4(_03597_),
    .ZN(_04743_));
 AOI221_X2 _21735_ (.A(_04741_),
    .B1(_04742_),
    .B2(net148),
    .C1(net86),
    .C2(_04743_),
    .ZN(_04744_));
 NAND3_X2 _21736_ (.A1(_04734_),
    .A2(_04739_),
    .A3(_04744_),
    .ZN(_04745_));
 NOR2_X1 _21737_ (.A1(_03530_),
    .A2(_03499_),
    .ZN(_04746_));
 NOR3_X4 _21738_ (.A1(_03510_),
    .A2(_04746_),
    .A3(_04737_),
    .ZN(_04747_));
 NOR2_X2 _21739_ (.A1(_04735_),
    .A2(_04737_),
    .ZN(_04748_));
 NOR2_X2 _21740_ (.A1(_03498_),
    .A2(_04245_),
    .ZN(_04749_));
 AOI222_X2 _21741_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_04747_),
    .B1(_04748_),
    .B2(\cs_registers_i.csr_mepc_o[23] ),
    .C1(_04749_),
    .C2(\cs_registers_i.dscratch1_q[23] ),
    .ZN(_04750_));
 CLKBUF_X2 _21742_ (.A(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .Z(_04751_));
 BUF_X4 _21743_ (.A(_04549_),
    .Z(_04752_));
 BUF_X4 _21744_ (.A(_04552_),
    .Z(_04753_));
 BUF_X2 _21745_ (.A(\cs_registers_i.mhpmcounter[2][55] ),
    .Z(_04754_));
 AOI22_X2 _21746_ (.A1(_04751_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04754_),
    .ZN(_04755_));
 OR2_X2 _21747_ (.A1(_03551_),
    .A2(_03536_),
    .ZN(_04756_));
 OAI21_X1 _21748_ (.A(_04750_),
    .B1(_04755_),
    .B2(_04756_),
    .ZN(_04757_));
 BUF_X2 _21749_ (.A(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .Z(_04758_));
 BUF_X2 _21750_ (.A(\cs_registers_i.mhpmcounter[2][23] ),
    .Z(_04759_));
 AOI22_X2 _21751_ (.A1(_04758_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04759_),
    .ZN(_04760_));
 NOR2_X1 _21752_ (.A1(_03532_),
    .A2(_04760_),
    .ZN(_04761_));
 OR3_X4 _21753_ (.A1(_04745_),
    .A2(_04757_),
    .A3(_04761_),
    .ZN(_04762_));
 OAI22_X4 _21754_ (.A1(_04661_),
    .A2(_04726_),
    .B1(_04762_),
    .B2(_04563_),
    .ZN(_04763_));
 BUF_X8 _21755_ (.A(_04263_),
    .Z(_04764_));
 AOI21_X4 _21756_ (.A(_04621_),
    .B1(_04763_),
    .B2(_04764_),
    .ZN(_04765_));
 BUF_X2 _21757_ (.A(_04765_),
    .Z(_04766_));
 MUX2_X1 _21758_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .S(_04615_),
    .Z(_01186_));
 MUX2_X1 _21759_ (.A(net40),
    .B(net48),
    .S(_04584_),
    .Z(_04767_));
 MUX2_X1 _21760_ (.A(net56),
    .B(net62),
    .S(_04584_),
    .Z(_04768_));
 MUX2_X1 _21761_ (.A(_04767_),
    .B(_04768_),
    .S(_04577_),
    .Z(_04769_));
 AOI21_X2 _21762_ (.A(_04580_),
    .B1(_04581_),
    .B2(_04769_),
    .ZN(_04770_));
 BUF_X4 _21763_ (.A(_04510_),
    .Z(_04771_));
 AOI211_X2 _21764_ (.A(_03502_),
    .B(_04509_),
    .C1(_03540_),
    .C2(_10922_),
    .ZN(_04772_));
 BUF_X4 _21765_ (.A(_04772_),
    .Z(_04773_));
 AOI22_X1 _21766_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_04771_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .ZN(_04774_));
 BUF_X4 _21767_ (.A(_04529_),
    .Z(_04775_));
 AOI22_X1 _21768_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(_04514_),
    .B1(_04775_),
    .B2(\cs_registers_i.dscratch1_q[27] ),
    .ZN(_04776_));
 AOI222_X2 _21769_ (.A1(net138),
    .A2(_04517_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[27] ),
    .C1(\cs_registers_i.mscratch_q[27] ),
    .C2(_04523_),
    .ZN(_04777_));
 OAI21_X1 _21770_ (.A(_04533_),
    .B1(_04536_),
    .B2(_00007_),
    .ZN(_04778_));
 AOI221_X2 _21771_ (.A(_04778_),
    .B1(_04526_),
    .B2(net90),
    .C1(\cs_registers_i.csr_mepc_o[27] ),
    .C2(_04543_),
    .ZN(_04779_));
 AND4_X1 _21772_ (.A1(_04774_),
    .A2(_04776_),
    .A3(_04777_),
    .A4(_04779_),
    .ZN(_04780_));
 BUF_X2 _21773_ (.A(\cs_registers_i.mhpmcounter[2][59] ),
    .Z(_04781_));
 AOI22_X4 _21774_ (.A1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(_04781_),
    .ZN(_04782_));
 BUF_X4 _21775_ (.A(_04559_),
    .Z(_04783_));
 BUF_X4 _21776_ (.A(_04752_),
    .Z(_04784_));
 BUF_X4 _21777_ (.A(_04753_),
    .Z(_04785_));
 AOI22_X2 _21778_ (.A1(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][27] ),
    .ZN(_04786_));
 OAI221_X2 _21779_ (.A(_04780_),
    .B1(_04782_),
    .B2(_04557_),
    .C1(_04783_),
    .C2(_04786_),
    .ZN(_04787_));
 NOR2_X1 _21780_ (.A1(_04393_),
    .A2(_04787_),
    .ZN(_04788_));
 MUX2_X2 _21781_ (.A(_04770_),
    .B(_04788_),
    .S(_04263_),
    .Z(_04789_));
 AOI21_X1 _21782_ (.A(_11408_),
    .B1(_03824_),
    .B2(net300),
    .ZN(_04790_));
 BUF_X4 _21783_ (.A(_04502_),
    .Z(_04791_));
 INV_X1 _21784_ (.A(_15793_),
    .ZN(_04792_));
 BUF_X1 _21785_ (.A(_15787_),
    .Z(_04793_));
 AOI21_X1 _21786_ (.A(_15786_),
    .B1(_15780_),
    .B2(_04793_),
    .ZN(_04794_));
 OR2_X1 _21787_ (.A1(_04792_),
    .A2(_04794_),
    .ZN(_04795_));
 NAND3_X2 _21788_ (.A1(_15781_),
    .A2(_04793_),
    .A3(_15793_),
    .ZN(_04796_));
 INV_X1 _21789_ (.A(_15774_),
    .ZN(_04797_));
 OAI21_X1 _21790_ (.A(_15775_),
    .B1(_15768_),
    .B2(_15769_),
    .ZN(_04798_));
 NAND2_X1 _21791_ (.A1(_04797_),
    .A2(_04798_),
    .ZN(_04799_));
 OR3_X1 _21792_ (.A1(_15762_),
    .A2(_15768_),
    .A3(_15774_),
    .ZN(_04800_));
 OAI21_X4 _21793_ (.A(_04799_),
    .B1(_04655_),
    .B2(_04800_),
    .ZN(_04801_));
 OAI21_X4 _21794_ (.A(_04795_),
    .B1(_04801_),
    .B2(_04796_),
    .ZN(_04802_));
 OAI21_X1 _21795_ (.A(_15799_),
    .B1(_15792_),
    .B2(_04802_),
    .ZN(_04803_));
 OR3_X4 _21796_ (.A1(_15799_),
    .A2(_04802_),
    .A3(_15792_),
    .ZN(_04804_));
 NAND3_X4 _21797_ (.A1(_04791_),
    .A2(_04803_),
    .A3(_04804_),
    .ZN(_04805_));
 INV_X1 _21798_ (.A(_04481_),
    .ZN(_04806_));
 INV_X1 _21799_ (.A(_15658_),
    .ZN(_04807_));
 NOR4_X2 _21800_ (.A1(_04806_),
    .A2(_04807_),
    .A3(_04646_),
    .A4(_04650_),
    .ZN(_04808_));
 NOR3_X2 _21801_ (.A1(_15671_),
    .A2(_04648_),
    .A3(_04808_),
    .ZN(_04809_));
 XNOR2_X2 _21802_ (.A(_04484_),
    .B(_04809_),
    .ZN(_04810_));
 OAI21_X4 _21803_ (.A(_04805_),
    .B1(_04810_),
    .B2(_04791_),
    .ZN(_04811_));
 OAI21_X4 _21804_ (.A(_04790_),
    .B1(_04811_),
    .B2(net300),
    .ZN(_04812_));
 AND4_X4 _21805_ (.A1(_04812_),
    .A2(_03439_),
    .A3(_04232_),
    .A4(_04563_),
    .ZN(_04813_));
 AND2_X1 _21806_ (.A1(_11406_),
    .A2(_04388_),
    .ZN(_04814_));
 BUF_X4 _21807_ (.A(_04814_),
    .Z(_04815_));
 OR2_X1 _21808_ (.A1(_04306_),
    .A2(_04685_),
    .ZN(_04816_));
 AND2_X1 _21809_ (.A1(_04275_),
    .A2(_04816_),
    .ZN(_04817_));
 OAI21_X1 _21810_ (.A(_15841_),
    .B1(_04297_),
    .B2(_04296_),
    .ZN(_04818_));
 OAI21_X1 _21811_ (.A(_10739_),
    .B1(_04297_),
    .B2(_04296_),
    .ZN(_04819_));
 OAI222_X2 _21812_ (.A1(_04409_),
    .A2(_04676_),
    .B1(_04818_),
    .B2(_04681_),
    .C1(_04819_),
    .C2(_04679_),
    .ZN(_04820_));
 NAND2_X1 _21813_ (.A1(_04685_),
    .A2(_04820_),
    .ZN(_04821_));
 NAND2_X1 _21814_ (.A1(_04817_),
    .A2(_04821_),
    .ZN(_04822_));
 AOI221_X1 _21815_ (.A(_04353_),
    .B1(_04360_),
    .B2(_16055_),
    .C1(_04363_),
    .C2(_16054_),
    .ZN(_04823_));
 AOI21_X1 _21816_ (.A(_04823_),
    .B1(_04370_),
    .B2(_16058_),
    .ZN(_04824_));
 BUF_X4 _21817_ (.A(_04368_),
    .Z(_04825_));
 AOI21_X1 _21818_ (.A(_04824_),
    .B1(_04825_),
    .B2(\alu_adder_result_ex[27] ),
    .ZN(_04826_));
 NAND2_X1 _21819_ (.A1(_04822_),
    .A2(_04826_),
    .ZN(_04827_));
 AOI21_X2 _21820_ (.A(_04408_),
    .B1(_04330_),
    .B2(_04693_),
    .ZN(_04828_));
 AOI221_X2 _21821_ (.A(_04292_),
    .B1(_04692_),
    .B2(_04828_),
    .C1(_04699_),
    .C2(_04409_),
    .ZN(_04829_));
 AOI21_X4 _21822_ (.A(_04673_),
    .B1(_04691_),
    .B2(_04410_),
    .ZN(_04830_));
 AOI21_X2 _21823_ (.A(_04829_),
    .B1(_04830_),
    .B2(_04292_),
    .ZN(_04831_));
 NAND3_X1 _21824_ (.A1(_04332_),
    .A2(_04702_),
    .A3(_04704_),
    .ZN(_04832_));
 OAI21_X1 _21825_ (.A(_04832_),
    .B1(_04711_),
    .B2(_04333_),
    .ZN(_04833_));
 NAND2_X1 _21826_ (.A1(_04332_),
    .A2(_04717_),
    .ZN(_04834_));
 MUX2_X1 _21827_ (.A(_15897_),
    .B(_16029_),
    .S(_04434_),
    .Z(_04835_));
 MUX2_X1 _21828_ (.A(_15889_),
    .B(_16040_),
    .S(_04434_),
    .Z(_04836_));
 MUX2_X1 _21829_ (.A(_04835_),
    .B(_04836_),
    .S(_10739_),
    .Z(_04837_));
 MUX2_X1 _21830_ (.A(_15881_),
    .B(_16045_),
    .S(_04434_),
    .Z(_04838_));
 NOR2_X1 _21831_ (.A1(_04397_),
    .A2(_04838_),
    .ZN(_04839_));
 CLKBUF_X3 _21832_ (.A(_04434_),
    .Z(_04840_));
 MUX2_X1 _21833_ (.A(_15868_),
    .B(_16052_),
    .S(_04840_),
    .Z(_04841_));
 AOI21_X1 _21834_ (.A(_04839_),
    .B1(_04841_),
    .B2(_04397_),
    .ZN(_04842_));
 MUX2_X1 _21835_ (.A(_04837_),
    .B(_04842_),
    .S(_04406_),
    .Z(_04843_));
 OAI22_X1 _21836_ (.A1(_04715_),
    .A2(_04834_),
    .B1(_04843_),
    .B2(_04333_),
    .ZN(_04844_));
 MUX2_X1 _21837_ (.A(_04833_),
    .B(_04844_),
    .S(_04452_),
    .Z(_04845_));
 MUX2_X1 _21838_ (.A(_04831_),
    .B(_04845_),
    .S(_04412_),
    .Z(_04846_));
 AND2_X1 _21839_ (.A1(_04457_),
    .A2(_04846_),
    .ZN(_04847_));
 OAI21_X2 _21840_ (.A(_04815_),
    .B1(_04827_),
    .B2(_04847_),
    .ZN(_04848_));
 AOI21_X4 _21841_ (.A(_04789_),
    .B1(_04813_),
    .B2(_04848_),
    .ZN(_04849_));
 BUF_X4 _21842_ (.A(_04849_),
    .Z(_04850_));
 NAND2_X2 _21843_ (.A1(_10394_),
    .A2(_10902_),
    .ZN(_04851_));
 NOR2_X4 _21844_ (.A1(_10903_),
    .A2(_04851_),
    .ZN(_04852_));
 NAND2_X1 _21845_ (.A1(_10900_),
    .A2(_10901_),
    .ZN(_04853_));
 AOI21_X4 _21846_ (.A(_04853_),
    .B1(_04605_),
    .B2(_04611_),
    .ZN(_04854_));
 NAND2_X4 _21847_ (.A1(_04852_),
    .A2(_04854_),
    .ZN(_04855_));
 MUX2_X1 _21848_ (.A(net333),
    .B(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(_04855_),
    .Z(_01187_));
 BUF_X4 _21849_ (.A(_04614_),
    .Z(_04856_));
 NAND2_X1 _21850_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .A2(_04856_),
    .ZN(_04857_));
 OR2_X2 _21851_ (.A1(_04573_),
    .A2(_04565_),
    .ZN(_04858_));
 BUF_X4 _21852_ (.A(_04858_),
    .Z(_04859_));
 MUX2_X1 _21853_ (.A(net67),
    .B(net45),
    .S(_04585_),
    .Z(_04860_));
 NAND2_X1 _21854_ (.A1(_04597_),
    .A2(_04860_),
    .ZN(_04861_));
 MUX2_X1 _21855_ (.A(net53),
    .B(net38),
    .S(_04585_),
    .Z(_04862_));
 NAND2_X1 _21856_ (.A1(_04619_),
    .A2(_04862_),
    .ZN(_04863_));
 AOI21_X2 _21857_ (.A(_04859_),
    .B1(_04861_),
    .B2(_04863_),
    .ZN(_04864_));
 AOI221_X1 _21858_ (.A(_04351_),
    .B1(_04358_),
    .B2(_16031_),
    .C1(_04362_),
    .C2(_16034_),
    .ZN(_04865_));
 AOI21_X1 _21859_ (.A(_04865_),
    .B1(_04353_),
    .B2(_16030_),
    .ZN(_04866_));
 NAND2_X1 _21860_ (.A1(_04685_),
    .A2(_04695_),
    .ZN(_04867_));
 AOI221_X2 _21861_ (.A(_04866_),
    .B1(_04867_),
    .B2(_04817_),
    .C1(_04369_),
    .C2(\alu_adder_result_ex[24] ),
    .ZN(_04868_));
 NOR2_X1 _21862_ (.A1(_04391_),
    .A2(_04868_),
    .ZN(_04869_));
 MUX2_X1 _21863_ (.A(_04439_),
    .B(_04448_),
    .S(_04712_),
    .Z(_04870_));
 MUX2_X1 _21864_ (.A(_04442_),
    .B(_04444_),
    .S(_15835_),
    .Z(_04871_));
 MUX2_X1 _21865_ (.A(_04713_),
    .B(_04835_),
    .S(_15835_),
    .Z(_04872_));
 MUX2_X1 _21866_ (.A(_04871_),
    .B(_04872_),
    .S(_04712_),
    .Z(_04873_));
 MUX2_X1 _21867_ (.A(_04870_),
    .B(_04873_),
    .S(_04707_),
    .Z(_04874_));
 AOI21_X1 _21868_ (.A(_04293_),
    .B1(_04874_),
    .B2(_04722_),
    .ZN(_04875_));
 OAI21_X1 _21869_ (.A(_04875_),
    .B1(_04684_),
    .B2(_04722_),
    .ZN(_04876_));
 AOI21_X1 _21870_ (.A(_04720_),
    .B1(_04677_),
    .B2(_04282_),
    .ZN(_04877_));
 MUX2_X1 _21871_ (.A(_04325_),
    .B(_04415_),
    .S(_10739_),
    .Z(_04878_));
 MUX2_X1 _21872_ (.A(_04878_),
    .B(_04428_),
    .S(_04406_),
    .Z(_04879_));
 OR2_X1 _21873_ (.A1(_04431_),
    .A2(_04879_),
    .ZN(_04880_));
 OAI21_X1 _21874_ (.A(_04424_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04881_));
 OAI21_X1 _21875_ (.A(_04881_),
    .B1(_04436_),
    .B2(_04429_),
    .ZN(_04882_));
 OAI21_X1 _21876_ (.A(_04880_),
    .B1(_04882_),
    .B2(_04333_),
    .ZN(_04883_));
 OAI21_X1 _21877_ (.A(_04877_),
    .B1(_04883_),
    .B2(_04282_),
    .ZN(_04884_));
 AOI21_X1 _21878_ (.A(_04725_),
    .B1(_04876_),
    .B2(_04884_),
    .ZN(_04885_));
 XNOR2_X2 _21879_ (.A(_04481_),
    .B(_04480_),
    .ZN(_04886_));
 INV_X1 _21880_ (.A(_15781_),
    .ZN(_04887_));
 OAI21_X4 _21881_ (.A(_04799_),
    .B1(_04800_),
    .B2(_04499_),
    .ZN(_04888_));
 XNOR2_X2 _21882_ (.A(_04887_),
    .B(_04888_),
    .ZN(_04889_));
 MUX2_X1 _21883_ (.A(_04886_),
    .B(_04889_),
    .S(_04463_),
    .Z(_04890_));
 MUX2_X1 _21884_ (.A(_03817_),
    .B(_04890_),
    .S(_12102_),
    .Z(_04891_));
 NOR2_X2 _21885_ (.A1(_11408_),
    .A2(_04891_),
    .ZN(_04892_));
 AOI22_X1 _21886_ (.A1(\cs_registers_i.dscratch0_q[24] ),
    .A2(_04771_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .ZN(_04893_));
 AOI22_X1 _21887_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(_04514_),
    .B1(_04775_),
    .B2(\cs_registers_i.dscratch1_q[24] ),
    .ZN(_04894_));
 AOI222_X2 _21888_ (.A1(net149),
    .A2(_04517_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[24] ),
    .C1(\cs_registers_i.mscratch_q[24] ),
    .C2(_04523_),
    .ZN(_04895_));
 OAI21_X1 _21889_ (.A(_04533_),
    .B1(_04536_),
    .B2(_01181_),
    .ZN(_04896_));
 AOI221_X1 _21890_ (.A(_04896_),
    .B1(_04526_),
    .B2(net87),
    .C1(\cs_registers_i.csr_mepc_o[24] ),
    .C2(_04543_),
    .ZN(_04897_));
 AND4_X1 _21891_ (.A1(_04893_),
    .A2(_04894_),
    .A3(_04895_),
    .A4(_04897_),
    .ZN(_04898_));
 BUF_X2 _21892_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .Z(_04899_));
 AOI22_X4 _21893_ (.A1(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(_04899_),
    .ZN(_04900_));
 BUF_X2 _21894_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .Z(_04901_));
 AOI22_X2 _21895_ (.A1(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A2(_04784_),
    .B1(_04785_),
    .B2(_04901_),
    .ZN(_04902_));
 OAI221_X2 _21896_ (.A(_04898_),
    .B1(_04900_),
    .B2(_04557_),
    .C1(_04783_),
    .C2(_04902_),
    .ZN(_04903_));
 OR4_X4 _21897_ (.A1(_04892_),
    .A2(_04885_),
    .A3(_04869_),
    .A4(_04903_),
    .ZN(_04904_));
 NAND3_X4 _21898_ (.A1(_03439_),
    .A2(_04232_),
    .A3(_04261_),
    .ZN(_04905_));
 BUF_X8 _21899_ (.A(_04905_),
    .Z(_04906_));
 OAI22_X4 _21900_ (.A1(_04617_),
    .A2(_04864_),
    .B1(_04906_),
    .B2(_04904_),
    .ZN(_04907_));
 BUF_X8 _21901_ (.A(_04907_),
    .Z(_04908_));
 BUF_X4 _21902_ (.A(_04614_),
    .Z(_04909_));
 OAI21_X1 _21903_ (.A(_04857_),
    .B1(_04908_),
    .B2(_04909_),
    .ZN(_01188_));
 NAND2_X1 _21904_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .A2(_04856_),
    .ZN(_04910_));
 CLKBUF_X3 _21905_ (.A(_04584_),
    .Z(_04911_));
 MUX2_X1 _21906_ (.A(net68),
    .B(net46),
    .S(_04911_),
    .Z(_04912_));
 MUX2_X1 _21907_ (.A(net54),
    .B(net49),
    .S(_04911_),
    .Z(_04913_));
 MUX2_X1 _21908_ (.A(_04912_),
    .B(_04913_),
    .S(_04619_),
    .Z(_04914_));
 AOI21_X1 _21909_ (.A(_04580_),
    .B1(_04583_),
    .B2(_04914_),
    .ZN(_04915_));
 NAND3_X1 _21910_ (.A1(_04316_),
    .A2(_04295_),
    .A3(_04703_),
    .ZN(_04916_));
 OAI21_X1 _21911_ (.A(_04697_),
    .B1(_04320_),
    .B2(_04318_),
    .ZN(_04917_));
 NAND2_X1 _21912_ (.A1(_04916_),
    .A2(_04917_),
    .ZN(_04918_));
 AND3_X1 _21913_ (.A1(_04316_),
    .A2(_04294_),
    .A3(_04710_),
    .ZN(_04919_));
 NAND2_X1 _21914_ (.A1(_10738_),
    .A2(_04423_),
    .ZN(_04920_));
 NAND2_X1 _21915_ (.A1(_10739_),
    .A2(_04700_),
    .ZN(_04921_));
 AOI22_X1 _21916_ (.A1(_04316_),
    .A2(_04295_),
    .B1(_04920_),
    .B2(_04921_),
    .ZN(_04922_));
 OR2_X1 _21917_ (.A1(_04919_),
    .A2(_04922_),
    .ZN(_04923_));
 MUX2_X1 _21918_ (.A(_04918_),
    .B(_04923_),
    .S(_04707_),
    .Z(_04924_));
 NAND2_X1 _21919_ (.A1(_04723_),
    .A2(_04924_),
    .ZN(_04925_));
 AOI21_X1 _21920_ (.A(_04672_),
    .B1(_04712_),
    .B2(_04707_),
    .ZN(_04926_));
 AOI211_X2 _21921_ (.A(_10738_),
    .B(_04341_),
    .C1(_04313_),
    .C2(_16080_),
    .ZN(_04927_));
 AOI21_X2 _21922_ (.A(_04927_),
    .B1(_04303_),
    .B2(_10738_),
    .ZN(_04928_));
 NOR2_X1 _21923_ (.A1(_04298_),
    .A2(_04928_),
    .ZN(_04929_));
 NOR3_X1 _21924_ (.A1(_04722_),
    .A2(_04926_),
    .A3(_04929_),
    .ZN(_04930_));
 NOR2_X2 _21925_ (.A1(_04720_),
    .A2(_04930_),
    .ZN(_04931_));
 OR2_X1 _21926_ (.A1(_04722_),
    .A2(_04340_),
    .ZN(_04932_));
 MUX2_X1 _21927_ (.A(_04714_),
    .B(_04837_),
    .S(_04712_),
    .Z(_04933_));
 OR2_X1 _21928_ (.A1(_04333_),
    .A2(_04933_),
    .ZN(_04934_));
 AND3_X1 _21929_ (.A1(_04316_),
    .A2(_04295_),
    .A3(_04716_),
    .ZN(_04935_));
 AOI21_X1 _21930_ (.A(_04935_),
    .B1(_04708_),
    .B2(_04330_),
    .ZN(_04936_));
 AOI21_X1 _21931_ (.A(_04282_),
    .B1(_04333_),
    .B2(_04936_),
    .ZN(_04937_));
 AOI21_X2 _21932_ (.A(_04293_),
    .B1(_04934_),
    .B2(_04937_),
    .ZN(_04938_));
 AOI22_X4 _21933_ (.A1(_04925_),
    .A2(_04931_),
    .B1(_04932_),
    .B2(_04938_),
    .ZN(_04939_));
 NOR2_X2 _21934_ (.A1(_04342_),
    .A2(_04939_),
    .ZN(_04940_));
 NOR2_X1 _21935_ (.A1(_04806_),
    .A2(_04650_),
    .ZN(_04941_));
 NOR2_X1 _21936_ (.A1(_15643_),
    .A2(_04941_),
    .ZN(_04942_));
 XNOR2_X2 _21937_ (.A(_04807_),
    .B(_04942_),
    .ZN(_04943_));
 NOR2_X1 _21938_ (.A1(_04502_),
    .A2(_04943_),
    .ZN(_04944_));
 NOR2_X1 _21939_ (.A1(_04622_),
    .A2(_04944_),
    .ZN(_04945_));
 INV_X1 _21940_ (.A(_15780_),
    .ZN(_04946_));
 OAI21_X4 _21941_ (.A(_04946_),
    .B1(_04801_),
    .B2(_04887_),
    .ZN(_04947_));
 XNOR2_X2 _21942_ (.A(_04947_),
    .B(_04793_),
    .ZN(_04948_));
 OAI21_X4 _21943_ (.A(_04945_),
    .B1(_04626_),
    .B2(_04948_),
    .ZN(_04949_));
 AOI21_X1 _21944_ (.A(_11407_),
    .B1(_03819_),
    .B2(net304),
    .ZN(_04950_));
 AOI21_X4 _21945_ (.A(_04662_),
    .B1(_04950_),
    .B2(_04949_),
    .ZN(_04951_));
 AND2_X1 _21946_ (.A1(_04685_),
    .A2(_04411_),
    .ZN(_04952_));
 NAND2_X1 _21947_ (.A1(_04276_),
    .A2(_04816_),
    .ZN(_04953_));
 AOI22_X1 _21948_ (.A1(_16039_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_16038_),
    .ZN(_04954_));
 NOR2_X1 _21949_ (.A1(_04370_),
    .A2(_04954_),
    .ZN(_04955_));
 INV_X1 _21950_ (.A(_16042_),
    .ZN(_04956_));
 AOI221_X2 _21951_ (.A(_04955_),
    .B1(_04369_),
    .B2(\alu_adder_result_ex[25] ),
    .C1(_04956_),
    .C2(_04370_),
    .ZN(_04957_));
 OAI221_X2 _21952_ (.A(_04951_),
    .B1(_04952_),
    .B2(_04953_),
    .C1(_04391_),
    .C2(_04957_),
    .ZN(_04958_));
 BUF_X8 _21953_ (.A(_04550_),
    .Z(_04959_));
 BUF_X4 _21954_ (.A(_04553_),
    .Z(_04960_));
 AOI22_X4 _21955_ (.A1(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][57] ),
    .ZN(_04961_));
 NOR2_X2 _21956_ (.A1(_04558_),
    .A2(_04961_),
    .ZN(_04962_));
 BUF_X4 _21957_ (.A(_04752_),
    .Z(_04963_));
 BUF_X4 _21958_ (.A(_04753_),
    .Z(_04964_));
 AOI22_X2 _21959_ (.A1(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][25] ),
    .ZN(_04965_));
 NOR2_X2 _21960_ (.A1(_04783_),
    .A2(_04965_),
    .ZN(_04966_));
 AOI222_X2 _21961_ (.A1(net150),
    .A2(_04518_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[25] ),
    .C1(_04544_),
    .C2(\cs_registers_i.csr_mepc_o[25] ),
    .ZN(_04967_));
 BUF_X4 _21962_ (.A(_04773_),
    .Z(_04968_));
 AOI22_X2 _21963_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(_04511_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .ZN(_04969_));
 AOI22_X4 _21964_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(_04515_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[25] ),
    .ZN(_04970_));
 OAI21_X1 _21965_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01182_),
    .ZN(_04971_));
 BUF_X4 _21966_ (.A(_04523_),
    .Z(_04972_));
 AOI221_X2 _21967_ (.A(_04971_),
    .B1(_04527_),
    .B2(net88),
    .C1(\cs_registers_i.mscratch_q[25] ),
    .C2(_04972_),
    .ZN(_04973_));
 NAND4_X4 _21968_ (.A1(_04967_),
    .A2(_04969_),
    .A3(_04970_),
    .A4(_04973_),
    .ZN(_04974_));
 OR3_X2 _21969_ (.A1(_04962_),
    .A2(_04966_),
    .A3(_04974_),
    .ZN(_04975_));
 OAI22_X4 _21970_ (.A1(_04958_),
    .A2(_04940_),
    .B1(_04975_),
    .B2(_04563_),
    .ZN(_04976_));
 MUX2_X2 _21971_ (.A(_04915_),
    .B(_04976_),
    .S(_04600_),
    .Z(_04977_));
 BUF_X8 _21972_ (.A(_04977_),
    .Z(_04978_));
 OAI21_X4 _21973_ (.A(_04910_),
    .B1(net442),
    .B2(_04909_),
    .ZN(_01189_));
 MUX2_X1 _21974_ (.A(net39),
    .B(net47),
    .S(_04911_),
    .Z(_04979_));
 MUX2_X1 _21975_ (.A(net55),
    .B(net59),
    .S(_04911_),
    .Z(_04980_));
 MUX2_X1 _21976_ (.A(_04979_),
    .B(_04980_),
    .S(_04619_),
    .Z(_04981_));
 AOI21_X2 _21977_ (.A(_04617_),
    .B1(_04981_),
    .B2(_04583_),
    .ZN(_04982_));
 BUF_X4 _21978_ (.A(_04362_),
    .Z(_04983_));
 AOI221_X1 _21979_ (.A(_04352_),
    .B1(_04359_),
    .B2(_16047_),
    .C1(_04983_),
    .C2(_16050_),
    .ZN(_04984_));
 AOI21_X1 _21980_ (.A(_04984_),
    .B1(_04370_),
    .B2(_16046_),
    .ZN(_04985_));
 AOI21_X1 _21981_ (.A(_04985_),
    .B1(_04825_),
    .B2(net384),
    .ZN(_04986_));
 NAND2_X2 _21982_ (.A1(_04412_),
    .A2(_04452_),
    .ZN(_04987_));
 OAI33_X1 _21983_ (.A1(_04322_),
    .A2(_04317_),
    .A3(_04818_),
    .B1(_04819_),
    .B2(_04335_),
    .B3(_04337_),
    .ZN(_04988_));
 MUX2_X1 _21984_ (.A(_04928_),
    .B(_04674_),
    .S(_04330_),
    .Z(_04989_));
 AOI21_X2 _21985_ (.A(_04988_),
    .B1(_04989_),
    .B2(_04332_),
    .ZN(_04990_));
 NOR2_X1 _21986_ (.A1(_04987_),
    .A2(_04990_),
    .ZN(_04991_));
 OAI21_X1 _21987_ (.A(_04986_),
    .B1(_04991_),
    .B2(_04953_),
    .ZN(_04992_));
 AND2_X1 _21988_ (.A1(_04815_),
    .A2(_04992_),
    .ZN(_04993_));
 INV_X1 _21989_ (.A(_15657_),
    .ZN(_04994_));
 AOI21_X1 _21990_ (.A(_15643_),
    .B1(_04480_),
    .B2(_04481_),
    .ZN(_04995_));
 OAI21_X1 _21991_ (.A(_04994_),
    .B1(_04995_),
    .B2(_04807_),
    .ZN(_04996_));
 XNOR2_X2 _21992_ (.A(_04486_),
    .B(_04996_),
    .ZN(_04997_));
 NOR2_X1 _21993_ (.A1(_04502_),
    .A2(_04997_),
    .ZN(_04998_));
 OAI21_X4 _21994_ (.A(_04946_),
    .B1(_04888_),
    .B2(_04887_),
    .ZN(_04999_));
 AOI21_X4 _21995_ (.A(_15786_),
    .B1(_04999_),
    .B2(_04793_),
    .ZN(_05000_));
 XNOR2_X2 _21996_ (.A(_15793_),
    .B(_05000_),
    .ZN(_05001_));
 AOI21_X2 _21997_ (.A(_04998_),
    .B1(_05001_),
    .B2(_04502_),
    .ZN(_05002_));
 MUX2_X1 _21998_ (.A(_01000_),
    .B(_05002_),
    .S(_12103_),
    .Z(_05003_));
 NOR2_X4 _21999_ (.A1(_11408_),
    .A2(_05003_),
    .ZN(_05004_));
 AND3_X1 _22000_ (.A1(_15841_),
    .A2(_04394_),
    .A3(_04395_),
    .ZN(_05005_));
 NAND3_X2 _22001_ (.A1(_04409_),
    .A2(_04398_),
    .A3(_04400_),
    .ZN(_05006_));
 OAI22_X4 _22002_ (.A1(_04409_),
    .A2(_04674_),
    .B1(_05005_),
    .B2(_05006_),
    .ZN(_05007_));
 MUX2_X1 _22003_ (.A(_04421_),
    .B(_04407_),
    .S(_04332_),
    .Z(_05008_));
 MUX2_X1 _22004_ (.A(_05007_),
    .B(_05008_),
    .S(_04452_),
    .Z(_05009_));
 MUX2_X1 _22005_ (.A(_04430_),
    .B(_04441_),
    .S(_04410_),
    .Z(_05010_));
 MUX2_X1 _22006_ (.A(_15901_),
    .B(_16020_),
    .S(_04434_),
    .Z(_05011_));
 MUX2_X1 _22007_ (.A(_15893_),
    .B(_16033_),
    .S(_04840_),
    .Z(_05012_));
 MUX2_X1 _22008_ (.A(_05011_),
    .B(_05012_),
    .S(_04397_),
    .Z(_05013_));
 OR2_X1 _22009_ (.A1(_15841_),
    .A2(_04838_),
    .ZN(_05014_));
 OAI21_X1 _22010_ (.A(_05014_),
    .B1(_04836_),
    .B2(_04397_),
    .ZN(_05015_));
 MUX2_X1 _22011_ (.A(_05013_),
    .B(_05015_),
    .S(_04712_),
    .Z(_05016_));
 MUX2_X1 _22012_ (.A(_04450_),
    .B(_05016_),
    .S(_04410_),
    .Z(_05017_));
 MUX2_X1 _22013_ (.A(_05010_),
    .B(_05017_),
    .S(_04453_),
    .Z(_05018_));
 MUX2_X1 _22014_ (.A(_05009_),
    .B(_05018_),
    .S(_04722_),
    .Z(_05019_));
 AND2_X1 _22015_ (.A1(_04457_),
    .A2(_05019_),
    .ZN(_05020_));
 AOI22_X1 _22016_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(_04511_),
    .B1(_04515_),
    .B2(\cs_registers_i.mie_q[10] ),
    .ZN(_05021_));
 BUF_X4 _22017_ (.A(_04520_),
    .Z(_05022_));
 AOI222_X2 _22018_ (.A1(net137),
    .A2(_04518_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[26] ),
    .C1(\cs_registers_i.mscratch_q[26] ),
    .C2(_04972_),
    .ZN(_05023_));
 AOI22_X1 _22019_ (.A1(net89),
    .A2(_04528_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[26] ),
    .ZN(_05024_));
 INV_X1 _22020_ (.A(\cs_registers_i.csr_depc_o[26] ),
    .ZN(_05025_));
 OAI221_X1 _22021_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01183_),
    .C1(_04539_),
    .C2(_05025_),
    .ZN(_05026_));
 AOI21_X1 _22022_ (.A(_05026_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .ZN(_05027_));
 AND4_X1 _22023_ (.A1(_05021_),
    .A2(_05023_),
    .A3(_05024_),
    .A4(_05027_),
    .ZN(_05028_));
 BUF_X2 _22024_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .Z(_05029_));
 AOI22_X2 _22025_ (.A1(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(_05029_),
    .ZN(_05030_));
 BUF_X4 _22026_ (.A(_04557_),
    .Z(_05031_));
 BUF_X2 _22027_ (.A(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .Z(_05032_));
 AOI22_X2 _22028_ (.A1(_05032_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][26] ),
    .ZN(_05033_));
 OAI221_X2 _22029_ (.A(_05028_),
    .B1(_05030_),
    .B2(_05031_),
    .C1(_04560_),
    .C2(_05033_),
    .ZN(_05034_));
 NOR4_X4 _22030_ (.A1(_05004_),
    .A2(_04993_),
    .A3(_05020_),
    .A4(_05034_),
    .ZN(_05035_));
 AOI21_X4 _22031_ (.A(_04982_),
    .B1(_05035_),
    .B2(_04764_),
    .ZN(_05036_));
 BUF_X4 _22032_ (.A(_05036_),
    .Z(_05037_));
 MUX2_X1 _22033_ (.A(net418),
    .B(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .S(_04615_),
    .Z(_01190_));
 MUX2_X1 _22034_ (.A(net333),
    .B(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .S(_04615_),
    .Z(_01191_));
 MUX2_X1 _22035_ (.A(net41),
    .B(net50),
    .S(_04593_),
    .Z(_05038_));
 MUX2_X1 _22036_ (.A(net57),
    .B(net63),
    .S(_04593_),
    .Z(_05039_));
 MUX2_X1 _22037_ (.A(_05038_),
    .B(_05039_),
    .S(_04619_),
    .Z(_05040_));
 AOI21_X2 _22038_ (.A(_04617_),
    .B1(_05040_),
    .B2(_04583_),
    .ZN(_05041_));
 NOR2_X1 _22039_ (.A1(_04707_),
    .A2(_04873_),
    .ZN(_05042_));
 MUX2_X1 _22040_ (.A(_15865_),
    .B(_16060_),
    .S(_04840_),
    .Z(_05043_));
 MUX2_X1 _22041_ (.A(_04841_),
    .B(_05043_),
    .S(_15835_),
    .Z(_05044_));
 NOR2_X1 _22042_ (.A1(_04429_),
    .A2(_05044_),
    .ZN(_05045_));
 NOR2_X1 _22043_ (.A1(_04712_),
    .A2(_05015_),
    .ZN(_05046_));
 NOR3_X1 _22044_ (.A1(_04333_),
    .A2(_05045_),
    .A3(_05046_),
    .ZN(_05047_));
 NOR3_X1 _22045_ (.A1(_04987_),
    .A2(_05042_),
    .A3(_05047_),
    .ZN(_05048_));
 MUX2_X1 _22046_ (.A(_04882_),
    .B(_04870_),
    .S(_04410_),
    .Z(_05049_));
 INV_X1 _22047_ (.A(_04670_),
    .ZN(_05050_));
 MUX2_X1 _22048_ (.A(_04324_),
    .B(_04328_),
    .S(_15841_),
    .Z(_05051_));
 MUX2_X1 _22049_ (.A(_04334_),
    .B(_04327_),
    .S(_10739_),
    .Z(_05052_));
 MUX2_X1 _22050_ (.A(_05051_),
    .B(_05052_),
    .S(_04330_),
    .Z(_05053_));
 MUX2_X1 _22051_ (.A(_05053_),
    .B(_04879_),
    .S(_04409_),
    .Z(_05054_));
 MUX2_X2 _22052_ (.A(_04820_),
    .B(_05054_),
    .S(_04452_),
    .Z(_05055_));
 AOI221_X2 _22053_ (.A(_05048_),
    .B1(_05049_),
    .B2(_05050_),
    .C1(_04282_),
    .C2(_05055_),
    .ZN(_05056_));
 NAND2_X1 _22054_ (.A1(_04457_),
    .A2(_05056_),
    .ZN(_05057_));
 AOI21_X1 _22055_ (.A(_04953_),
    .B1(_04830_),
    .B2(_04685_),
    .ZN(_05058_));
 AOI221_X1 _22056_ (.A(_04352_),
    .B1(_04359_),
    .B2(_16063_),
    .C1(_04983_),
    .C2(_16062_),
    .ZN(_05059_));
 AOI21_X1 _22057_ (.A(_05059_),
    .B1(_04370_),
    .B2(_16066_),
    .ZN(_05060_));
 AOI21_X1 _22058_ (.A(_05060_),
    .B1(_04825_),
    .B2(\alu_adder_result_ex[28] ),
    .ZN(_05061_));
 INV_X1 _22059_ (.A(_05061_),
    .ZN(_05062_));
 OAI21_X1 _22060_ (.A(_04815_),
    .B1(_05058_),
    .B2(_05062_),
    .ZN(_05063_));
 AOI22_X2 _22061_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][60] ),
    .ZN(_05064_));
 NOR2_X1 _22062_ (.A1(_05031_),
    .A2(_05064_),
    .ZN(_05065_));
 BUF_X2 _22063_ (.A(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .Z(_05066_));
 BUF_X2 _22064_ (.A(\cs_registers_i.mhpmcounter[2][28] ),
    .Z(_05067_));
 AOI22_X1 _22065_ (.A1(_05066_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(_05067_),
    .ZN(_05068_));
 NOR2_X1 _22066_ (.A1(_04783_),
    .A2(_05068_),
    .ZN(_05069_));
 AOI22_X2 _22067_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(_04511_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .ZN(_05070_));
 AOI22_X2 _22068_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(_04515_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[28] ),
    .ZN(_05071_));
 AOI222_X2 _22069_ (.A1(net139),
    .A2(_04518_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[28] ),
    .C1(\cs_registers_i.mscratch_q[28] ),
    .C2(_04972_),
    .ZN(_05072_));
 OAI21_X1 _22070_ (.A(_04533_),
    .B1(_04536_),
    .B2(_00008_),
    .ZN(_05073_));
 BUF_X4 _22071_ (.A(_04543_),
    .Z(_05074_));
 AOI221_X2 _22072_ (.A(_05073_),
    .B1(_04527_),
    .B2(net91),
    .C1(\cs_registers_i.csr_mepc_o[28] ),
    .C2(_05074_),
    .ZN(_05075_));
 NAND4_X4 _22073_ (.A1(_05070_),
    .A2(_05071_),
    .A3(_05072_),
    .A4(_05075_),
    .ZN(_05076_));
 NOR3_X4 _22074_ (.A1(_05065_),
    .A2(_05069_),
    .A3(_05076_),
    .ZN(_05077_));
 NAND2_X1 _22075_ (.A1(net300),
    .A2(_03827_),
    .ZN(_05078_));
 CLKBUF_X3 _22076_ (.A(_04625_),
    .Z(_05079_));
 NOR2_X1 _22077_ (.A1(_15685_),
    .A2(_04488_),
    .ZN(_05080_));
 NOR2_X1 _22078_ (.A1(_04482_),
    .A2(_05080_),
    .ZN(_05081_));
 XOR2_X2 _22079_ (.A(net328),
    .B(_05081_),
    .Z(_05082_));
 NAND2_X1 _22080_ (.A1(_05079_),
    .A2(_05082_),
    .ZN(_05083_));
 INV_X1 _22081_ (.A(_15792_),
    .ZN(_05084_));
 AND2_X1 _22082_ (.A1(_05084_),
    .A2(_04795_),
    .ZN(_05085_));
 OAI21_X2 _22083_ (.A(_05085_),
    .B1(_04888_),
    .B2(_04796_),
    .ZN(_05086_));
 AOI21_X2 _22084_ (.A(_15798_),
    .B1(_15799_),
    .B2(_05086_),
    .ZN(_05087_));
 XOR2_X1 _22085_ (.A(_05087_),
    .B(_15805_),
    .Z(_05088_));
 OAI21_X2 _22086_ (.A(_05083_),
    .B1(_05079_),
    .B2(_05088_),
    .ZN(_05089_));
 OAI21_X2 _22087_ (.A(_05078_),
    .B1(_04622_),
    .B2(_05089_),
    .ZN(_05090_));
 OR2_X4 _22088_ (.A1(_05090_),
    .A2(_11408_),
    .ZN(_05091_));
 AND4_X4 _22089_ (.A1(_05091_),
    .A2(_05063_),
    .A3(_05077_),
    .A4(_05057_),
    .ZN(_05092_));
 AOI21_X4 _22090_ (.A(_05041_),
    .B1(_04764_),
    .B2(_05092_),
    .ZN(_05093_));
 BUF_X4 _22091_ (.A(_05093_),
    .Z(_05094_));
 MUX2_X1 _22092_ (.A(_05094_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .S(_04615_),
    .Z(_01192_));
 NAND2_X1 _22093_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(_04856_),
    .ZN(_05095_));
 MUX2_X1 _22094_ (.A(net42),
    .B(net51),
    .S(_04585_),
    .Z(_05096_));
 MUX2_X1 _22095_ (.A(net58),
    .B(net64),
    .S(_04585_),
    .Z(_05097_));
 MUX2_X1 _22096_ (.A(_05096_),
    .B(_05097_),
    .S(_04619_),
    .Z(_05098_));
 AOI21_X1 _22097_ (.A(_04617_),
    .B1(_05098_),
    .B2(_04583_),
    .ZN(_05099_));
 NAND2_X1 _22098_ (.A1(net300),
    .A2(_01093_),
    .ZN(_05100_));
 INV_X1 _22099_ (.A(_15699_),
    .ZN(_05101_));
 OAI21_X2 _22100_ (.A(_15700_),
    .B1(_15685_),
    .B2(_04652_),
    .ZN(_05102_));
 NAND2_X2 _22101_ (.A1(_05102_),
    .A2(_05101_),
    .ZN(_05103_));
 XOR2_X2 _22102_ (.A(_04491_),
    .B(_05103_),
    .Z(_05104_));
 NOR3_X1 _22103_ (.A1(_15799_),
    .A2(_15798_),
    .A3(_15804_),
    .ZN(_05105_));
 NOR2_X1 _22104_ (.A1(_15805_),
    .A2(_15804_),
    .ZN(_05106_));
 NOR2_X2 _22105_ (.A1(_05105_),
    .A2(_05106_),
    .ZN(_05107_));
 OR3_X1 _22106_ (.A1(_15792_),
    .A2(_15798_),
    .A3(_15804_),
    .ZN(_05108_));
 OAI21_X4 _22107_ (.A(_05107_),
    .B1(_04802_),
    .B2(_05108_),
    .ZN(_05109_));
 XNOR2_X2 _22108_ (.A(_15811_),
    .B(_05109_),
    .ZN(_05110_));
 MUX2_X1 _22109_ (.A(_05104_),
    .B(_05110_),
    .S(_04502_),
    .Z(_05111_));
 OAI21_X4 _22110_ (.A(_05100_),
    .B1(_05111_),
    .B2(net300),
    .ZN(_05112_));
 NOR2_X4 _22111_ (.A1(_05112_),
    .A2(_11409_),
    .ZN(_05113_));
 AOI22_X1 _22112_ (.A1(_16071_),
    .A2(_04359_),
    .B1(_04362_),
    .B2(_16070_),
    .ZN(_05114_));
 MUX2_X1 _22113_ (.A(_16074_),
    .B(_05114_),
    .S(_04664_),
    .Z(_05115_));
 NAND3_X1 _22114_ (.A1(_04281_),
    .A2(_04307_),
    .A3(_04275_),
    .ZN(_05116_));
 NAND2_X1 _22115_ (.A1(net14),
    .A2(_04368_),
    .ZN(_05117_));
 NAND3_X1 _22116_ (.A1(_05115_),
    .A2(_05116_),
    .A3(_05117_),
    .ZN(_05118_));
 MUX2_X2 _22117_ (.A(_04307_),
    .B(_05007_),
    .S(_04452_),
    .Z(_05119_));
 NOR2_X4 _22118_ (.A1(_04282_),
    .A2(_04687_),
    .ZN(_05120_));
 AOI21_X2 _22119_ (.A(_05118_),
    .B1(_05119_),
    .B2(_05120_),
    .ZN(_05121_));
 MUX2_X1 _22120_ (.A(_04331_),
    .B(_04918_),
    .S(_04408_),
    .Z(_05122_));
 MUX2_X1 _22121_ (.A(_15861_),
    .B(_16064_),
    .S(_04434_),
    .Z(_05123_));
 MUX2_X1 _22122_ (.A(_15856_),
    .B(_16072_),
    .S(_04434_),
    .Z(_05124_));
 MUX2_X1 _22123_ (.A(_05123_),
    .B(_05124_),
    .S(_04397_),
    .Z(_05125_));
 MUX2_X1 _22124_ (.A(_04842_),
    .B(_05125_),
    .S(_04712_),
    .Z(_05126_));
 MUX2_X1 _22125_ (.A(_04933_),
    .B(_05126_),
    .S(_04410_),
    .Z(_05127_));
 AOI22_X2 _22126_ (.A1(_04413_),
    .A2(_05122_),
    .B1(_05127_),
    .B2(_04685_),
    .ZN(_05128_));
 NOR3_X1 _22127_ (.A1(_04409_),
    .A2(_04919_),
    .A3(_04922_),
    .ZN(_05129_));
 AOI21_X1 _22128_ (.A(_05129_),
    .B1(_04936_),
    .B2(_04409_),
    .ZN(_05130_));
 NAND3_X1 _22129_ (.A1(_04412_),
    .A2(_04293_),
    .A3(_05130_),
    .ZN(_05131_));
 OR3_X1 _22130_ (.A1(_04412_),
    .A2(_04452_),
    .A3(_04990_),
    .ZN(_05132_));
 NAND4_X2 _22131_ (.A1(_04456_),
    .A2(_05128_),
    .A3(_05131_),
    .A4(_05132_),
    .ZN(_05133_));
 AOI221_X2 _22132_ (.A(_04390_),
    .B1(_05121_),
    .B2(_05133_),
    .C1(_10742_),
    .C2(_10661_),
    .ZN(_05134_));
 AOI22_X1 _22133_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(_04515_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .ZN(_05135_));
 AOI222_X2 _22134_ (.A1(net140),
    .A2(_04518_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[29] ),
    .C1(_05074_),
    .C2(\cs_registers_i.csr_mepc_o[29] ),
    .ZN(_05136_));
 AOI22_X1 _22135_ (.A1(net92),
    .A2(_04528_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[29] ),
    .ZN(_05137_));
 OAI21_X1 _22136_ (.A(_04534_),
    .B1(_04537_),
    .B2(_00009_),
    .ZN(_05138_));
 AOI221_X1 _22137_ (.A(_05138_),
    .B1(_04523_),
    .B2(\cs_registers_i.mscratch_q[29] ),
    .C1(\cs_registers_i.dscratch0_q[29] ),
    .C2(_04771_),
    .ZN(_05139_));
 AND4_X1 _22138_ (.A1(_05135_),
    .A2(_05136_),
    .A3(_05137_),
    .A4(_05139_),
    .ZN(_05140_));
 AOI22_X2 _22139_ (.A1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][61] ),
    .ZN(_05141_));
 BUF_X2 _22140_ (.A(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .Z(_05142_));
 CLKBUF_X2 _22141_ (.A(\cs_registers_i.mhpmcounter[2][29] ),
    .Z(_05143_));
 AOI22_X2 _22142_ (.A1(_05142_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(_05143_),
    .ZN(_05144_));
 OAI221_X2 _22143_ (.A(_05140_),
    .B1(_05141_),
    .B2(_04558_),
    .C1(_04560_),
    .C2(_05144_),
    .ZN(_05145_));
 NOR4_X4 _22144_ (.A1(_05113_),
    .A2(_04906_),
    .A3(_05134_),
    .A4(_05145_),
    .ZN(_05146_));
 OR2_X4 _22145_ (.A1(_05146_),
    .A2(_05099_),
    .ZN(_05147_));
 BUF_X16 _22146_ (.A(_05147_),
    .Z(_05148_));
 OAI21_X4 _22147_ (.A(_05095_),
    .B1(net445),
    .B2(_04909_),
    .ZN(_01193_));
 NAND2_X1 _22148_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_04369_),
    .ZN(_05149_));
 AOI22_X1 _22149_ (.A1(_16079_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_16078_),
    .ZN(_05150_));
 MUX2_X1 _22150_ (.A(_16082_),
    .B(_05150_),
    .S(_04665_),
    .Z(_05151_));
 AOI221_X2 _22151_ (.A(_04298_),
    .B1(_04290_),
    .B2(_04284_),
    .C1(_04279_),
    .C2(_04280_),
    .ZN(_05152_));
 MUX2_X1 _22152_ (.A(_04674_),
    .B(_04928_),
    .S(_05152_),
    .Z(_05153_));
 OAI211_X2 _22153_ (.A(_05149_),
    .B(_05151_),
    .C1(_05153_),
    .C2(_04687_),
    .ZN(_05154_));
 AOI21_X4 _22154_ (.A(_11407_),
    .B1(_01124_),
    .B2(_04622_),
    .ZN(_05155_));
 OAI21_X1 _22155_ (.A(_05101_),
    .B1(_04482_),
    .B2(_04489_),
    .ZN(_05156_));
 AOI21_X2 _22156_ (.A(_15706_),
    .B1(_05156_),
    .B2(_04491_),
    .ZN(_05157_));
 XNOR2_X2 _22157_ (.A(_15717_),
    .B(_05157_),
    .ZN(_05158_));
 AND2_X1 _22158_ (.A1(_04625_),
    .A2(_05158_),
    .ZN(_05159_));
 INV_X1 _22159_ (.A(_05108_),
    .ZN(_05160_));
 OAI221_X2 _22160_ (.A(_05160_),
    .B1(_04888_),
    .B2(_04796_),
    .C1(_04792_),
    .C2(_04794_),
    .ZN(_05161_));
 INV_X1 _22161_ (.A(_15811_),
    .ZN(_05162_));
 CLKBUF_X2 _22162_ (.A(_15817_),
    .Z(_05163_));
 NOR3_X1 _22163_ (.A1(_05162_),
    .A2(_05163_),
    .A3(_04624_),
    .ZN(_05164_));
 AND3_X4 _22164_ (.A1(_05107_),
    .A2(_05164_),
    .A3(_05161_),
    .ZN(_05165_));
 INV_X1 _22165_ (.A(_15810_),
    .ZN(_05166_));
 NAND3_X1 _22166_ (.A1(_05163_),
    .A2(_05166_),
    .A3(_04463_),
    .ZN(_05167_));
 AOI21_X2 _22167_ (.A(_05167_),
    .B1(_05107_),
    .B2(_05161_),
    .ZN(_05168_));
 NAND3_X1 _22168_ (.A1(_05162_),
    .A2(_05163_),
    .A3(_05166_),
    .ZN(_05169_));
 INV_X1 _22169_ (.A(_05163_),
    .ZN(_05170_));
 NAND2_X1 _22170_ (.A1(_05170_),
    .A2(_15810_),
    .ZN(_05171_));
 AOI21_X2 _22171_ (.A(_04624_),
    .B1(_05169_),
    .B2(_05171_),
    .ZN(_05172_));
 NOR4_X4 _22172_ (.A1(_05159_),
    .A2(_05165_),
    .A3(_05168_),
    .A4(_05172_),
    .ZN(_05173_));
 NAND2_X2 _22173_ (.A1(_12103_),
    .A2(_05173_),
    .ZN(_05174_));
 AOI22_X4 _22174_ (.A1(_04815_),
    .A2(_05154_),
    .B1(_05155_),
    .B2(_05174_),
    .ZN(_05175_));
 AOI211_X2 _22175_ (.A(_04332_),
    .B(_04425_),
    .C1(_04428_),
    .C2(_04330_),
    .ZN(_05176_));
 AOI221_X2 _22176_ (.A(_05176_),
    .B1(_04290_),
    .B2(_04284_),
    .C1(_04332_),
    .C2(_04421_),
    .ZN(_05177_));
 AOI211_X2 _22177_ (.A(_04412_),
    .B(_05177_),
    .C1(_04411_),
    .C2(_04293_),
    .ZN(_05178_));
 MUX2_X1 _22178_ (.A(_15852_),
    .B(_16068_),
    .S(_04840_),
    .Z(_05179_));
 NAND2_X1 _22179_ (.A1(_15845_),
    .A2(_04342_),
    .ZN(_05180_));
 OAI21_X1 _22180_ (.A(_05180_),
    .B1(_04342_),
    .B2(_16080_),
    .ZN(_05181_));
 MUX2_X1 _22181_ (.A(_05179_),
    .B(_05181_),
    .S(_15835_),
    .Z(_05182_));
 MUX2_X1 _22182_ (.A(_05044_),
    .B(_05182_),
    .S(_04712_),
    .Z(_05183_));
 MUX2_X1 _22183_ (.A(_05016_),
    .B(_05183_),
    .S(_04707_),
    .Z(_05184_));
 MUX2_X1 _22184_ (.A(_04451_),
    .B(_05184_),
    .S(_04453_),
    .Z(_05185_));
 AOI21_X2 _22185_ (.A(_05178_),
    .B1(_05185_),
    .B2(_04723_),
    .ZN(_05186_));
 OAI221_X2 _22186_ (.A(_05175_),
    .B1(_05186_),
    .B2(_04342_),
    .C1(_03465_),
    .C2(_10678_),
    .ZN(_05187_));
 CLKBUF_X2 _22187_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .Z(_05188_));
 AOI22_X2 _22188_ (.A1(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(_05188_),
    .ZN(_05189_));
 NOR3_X2 _22189_ (.A1(_03551_),
    .A2(_04236_),
    .A3(_05189_),
    .ZN(_05190_));
 AOI22_X1 _22190_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(\cs_registers_i.mhpmcounter[2][30] ),
    .ZN(_05191_));
 NOR2_X1 _22191_ (.A1(_04559_),
    .A2(_05191_),
    .ZN(_05192_));
 AOI22_X2 _22192_ (.A1(net141),
    .A2(_04518_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[30] ),
    .ZN(_05193_));
 AOI22_X2 _22193_ (.A1(\cs_registers_i.mscratch_q[30] ),
    .A2(_04524_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[30] ),
    .ZN(_05194_));
 NAND2_X2 _22194_ (.A1(_05193_),
    .A2(_05194_),
    .ZN(_05195_));
 AOI22_X2 _22195_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(_04515_),
    .B1(_04775_),
    .B2(\cs_registers_i.dscratch1_q[30] ),
    .ZN(_05196_));
 AOI22_X2 _22196_ (.A1(net94),
    .A2(_04528_),
    .B1(_04771_),
    .B2(\cs_registers_i.dscratch0_q[30] ),
    .ZN(_05197_));
 AOI211_X2 _22197_ (.A(_03500_),
    .B(_04509_),
    .C1(_03518_),
    .C2(_03540_),
    .ZN(_05198_));
 AND4_X4 _22198_ (.A1(_11065_),
    .A2(_03594_),
    .A3(_04249_),
    .A4(_04535_),
    .ZN(_05199_));
 INV_X1 _22199_ (.A(_00010_),
    .ZN(_05200_));
 AOI221_X2 _22200_ (.A(net17),
    .B1(_05199_),
    .B2(_05200_),
    .C1(\cs_registers_i.csr_depc_o[30] ),
    .C2(_04772_),
    .ZN(_05201_));
 NAND4_X4 _22201_ (.A1(_04247_),
    .A2(_05196_),
    .A3(_05197_),
    .A4(_05201_),
    .ZN(_05202_));
 NOR4_X4 _22202_ (.A1(_05190_),
    .A2(_05192_),
    .A3(_05195_),
    .A4(_05202_),
    .ZN(_05203_));
 NAND2_X1 _22203_ (.A1(_04662_),
    .A2(_05203_),
    .ZN(_05204_));
 AOI21_X4 _22204_ (.A(_04906_),
    .B1(_05187_),
    .B2(_05204_),
    .ZN(_05205_));
 MUX2_X1 _22205_ (.A(net43),
    .B(net52),
    .S(_04584_),
    .Z(_05206_));
 MUX2_X1 _22206_ (.A(net60),
    .B(net65),
    .S(_04584_),
    .Z(_05207_));
 MUX2_X1 _22207_ (.A(_05206_),
    .B(_05207_),
    .S(_04619_),
    .Z(_05208_));
 AOI21_X4 _22208_ (.A(_04580_),
    .B1(_04583_),
    .B2(_05208_),
    .ZN(_05209_));
 AOI21_X4 _22209_ (.A(_05205_),
    .B1(_05209_),
    .B2(_04906_),
    .ZN(_05210_));
 BUF_X4 _22210_ (.A(_05210_),
    .Z(_05211_));
 MUX2_X1 _22211_ (.A(_05211_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .S(_04615_),
    .Z(_01194_));
 NAND2_X1 _22212_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(_04856_),
    .ZN(_05212_));
 NOR2_X1 _22213_ (.A1(_04597_),
    .A2(_04575_),
    .ZN(_05213_));
 NOR2_X1 _22214_ (.A1(_04619_),
    .A2(_04576_),
    .ZN(_05214_));
 NOR3_X2 _22215_ (.A1(_04859_),
    .A2(_05213_),
    .A3(_05214_),
    .ZN(_05215_));
 AOI21_X2 _22216_ (.A(_15706_),
    .B1(_05103_),
    .B2(_04491_),
    .ZN(_05216_));
 INV_X1 _22217_ (.A(_15717_),
    .ZN(_05217_));
 OAI21_X2 _22218_ (.A(_04639_),
    .B1(_05216_),
    .B2(_05217_),
    .ZN(_05218_));
 XNOR2_X2 _22219_ (.A(_15726_),
    .B(_05218_),
    .ZN(_05219_));
 OAI21_X1 _22220_ (.A(_12103_),
    .B1(_04791_),
    .B2(_05219_),
    .ZN(_05220_));
 OAI21_X4 _22221_ (.A(_05166_),
    .B1(_05109_),
    .B2(_05162_),
    .ZN(_05221_));
 AOI21_X4 _22222_ (.A(_15816_),
    .B1(_05221_),
    .B2(_05163_),
    .ZN(_05222_));
 XNOR2_X2 _22223_ (.A(_05222_),
    .B(_15823_),
    .ZN(_05223_));
 AOI21_X2 _22224_ (.A(_05220_),
    .B1(_05223_),
    .B2(_04791_),
    .ZN(_05224_));
 AND2_X1 _22225_ (.A1(net300),
    .A2(_03412_),
    .ZN(_05225_));
 NOR3_X4 _22226_ (.A1(_05225_),
    .A2(_11409_),
    .A3(_05224_),
    .ZN(_05226_));
 NAND2_X1 _22227_ (.A1(\cs_registers_i.csr_mepc_o[31] ),
    .A2(_04542_),
    .ZN(_05227_));
 AOI211_X2 _22228_ (.A(_03504_),
    .B(_04244_),
    .C1(_03518_),
    .C2(_03540_),
    .ZN(_05228_));
 AOI222_X2 _22229_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(_04519_),
    .B1(_05228_),
    .B2(\cs_registers_i.mcause_q[5] ),
    .C1(\cs_registers_i.mscratch_q[31] ),
    .C2(_04522_),
    .ZN(_05229_));
 AOI222_X2 _22230_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_04529_),
    .B1(_04772_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .C1(net95),
    .C2(_04526_),
    .ZN(_05230_));
 NOR3_X4 _22231_ (.A1(_03580_),
    .A2(_03581_),
    .A3(_04512_),
    .ZN(_05231_));
 INV_X1 _22232_ (.A(_00011_),
    .ZN(_05232_));
 AOI221_X1 _22233_ (.A(_05231_),
    .B1(_05199_),
    .B2(_05232_),
    .C1(net16),
    .C2(\cs_registers_i.dscratch0_q[31] ),
    .ZN(_05233_));
 AND4_X1 _22234_ (.A1(_05227_),
    .A2(_05229_),
    .A3(_05230_),
    .A4(_05233_),
    .ZN(_05234_));
 AOI22_X4 _22235_ (.A1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .A2(_04549_),
    .B1(_04552_),
    .B2(\cs_registers_i.mhpmcounter[2][63] ),
    .ZN(_05235_));
 BUF_X2 _22236_ (.A(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .Z(_05236_));
 AOI22_X2 _22237_ (.A1(_05236_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(\cs_registers_i.mhpmcounter[2][31] ),
    .ZN(_05237_));
 OAI221_X2 _22238_ (.A(_05234_),
    .B1(_05235_),
    .B2(_04556_),
    .C1(_04235_),
    .C2(_05237_),
    .ZN(_05238_));
 NAND2_X1 _22239_ (.A1(_04410_),
    .A2(_04685_),
    .ZN(_05239_));
 MUX2_X1 _22240_ (.A(_04676_),
    .B(_04306_),
    .S(_05239_),
    .Z(_05240_));
 CLKBUF_X3 _22241_ (.A(_15494_),
    .Z(_05241_));
 AOI221_X1 _22242_ (.A(_04350_),
    .B1(_04358_),
    .B2(_05241_),
    .C1(_04361_),
    .C2(_15497_),
    .ZN(_05242_));
 AOI21_X1 _22243_ (.A(_05242_),
    .B1(_04352_),
    .B2(_15493_),
    .ZN(_05243_));
 AND2_X1 _22244_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_04367_),
    .ZN(_05244_));
 OR2_X1 _22245_ (.A1(_05243_),
    .A2(_05244_),
    .ZN(_05245_));
 AOI221_X2 _22246_ (.A(_05238_),
    .B1(_05240_),
    .B2(_04276_),
    .C1(_04815_),
    .C2(_05245_),
    .ZN(_05246_));
 NAND2_X1 _22247_ (.A1(_04282_),
    .A2(_04453_),
    .ZN(_05247_));
 MUX2_X1 _22248_ (.A(_15842_),
    .B(_15496_),
    .S(_04840_),
    .Z(_05248_));
 MUX2_X1 _22249_ (.A(_05181_),
    .B(_05248_),
    .S(_15835_),
    .Z(_05249_));
 NAND3_X1 _22250_ (.A1(_04431_),
    .A2(_04712_),
    .A3(_05249_),
    .ZN(_05250_));
 NAND2_X1 _22251_ (.A1(_04431_),
    .A2(_04429_),
    .ZN(_05251_));
 OAI221_X1 _22252_ (.A(_05250_),
    .B1(_05251_),
    .B2(_05125_),
    .C1(_04843_),
    .C2(_04707_),
    .ZN(_05252_));
 OAI22_X1 _22253_ (.A1(_05247_),
    .A2(_04706_),
    .B1(_05252_),
    .B2(_04987_),
    .ZN(_05253_));
 NOR2_X1 _22254_ (.A1(_04670_),
    .A2(_04719_),
    .ZN(_05254_));
 AND3_X1 _22255_ (.A1(_04282_),
    .A2(_04293_),
    .A3(_04695_),
    .ZN(_05255_));
 OR3_X1 _22256_ (.A1(_05253_),
    .A2(_05254_),
    .A3(_05255_),
    .ZN(_05256_));
 OAI21_X2 _22257_ (.A(_05246_),
    .B1(_05256_),
    .B2(_04725_),
    .ZN(_05257_));
 OR2_X1 _22258_ (.A1(_04905_),
    .A2(_05257_),
    .ZN(_05258_));
 OAI22_X4 _22259_ (.A1(_04617_),
    .A2(_05215_),
    .B1(_05226_),
    .B2(_05258_),
    .ZN(_05259_));
 BUF_X8 _22260_ (.A(_05259_),
    .Z(_05260_));
 OAI21_X4 _22261_ (.A(_05212_),
    .B1(net441),
    .B2(_04909_),
    .ZN(_01195_));
 CLKBUF_X3 _22262_ (.A(_04589_),
    .Z(_05261_));
 NOR2_X4 _22263_ (.A1(_04570_),
    .A2(_04588_),
    .ZN(_05262_));
 AND2_X1 _22264_ (.A1(_04589_),
    .A2(net45),
    .ZN(_05263_));
 AOI221_X2 _22265_ (.A(_04581_),
    .B1(_05262_),
    .B2(net67),
    .C1(_05263_),
    .C2(_04570_),
    .ZN(_05264_));
 NOR2_X4 _22266_ (.A1(_04577_),
    .A2(_04584_),
    .ZN(_05265_));
 AOI221_X2 _22267_ (.A(_04858_),
    .B1(_05262_),
    .B2(\load_store_unit_i.rdata_q[8] ),
    .C1(_05265_),
    .C2(\load_store_unit_i.rdata_q[16] ),
    .ZN(_05266_));
 NOR3_X1 _22268_ (.A1(_05261_),
    .A2(_05264_),
    .A3(_05266_),
    .ZN(_05267_));
 CLKBUF_X3 _22269_ (.A(_04570_),
    .Z(_05268_));
 NOR2_X1 _22270_ (.A1(_05268_),
    .A2(_04586_),
    .ZN(_05269_));
 BUF_X4 _22271_ (.A(_04565_),
    .Z(_05270_));
 INV_X1 _22272_ (.A(_04573_),
    .ZN(_05271_));
 NAND2_X4 _22273_ (.A1(_05271_),
    .A2(_04565_),
    .ZN(_05272_));
 AOI22_X2 _22274_ (.A1(_05270_),
    .A2(net53),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[24] ),
    .ZN(_05273_));
 OAI22_X2 _22275_ (.A1(_05264_),
    .A2(_05266_),
    .B1(_05273_),
    .B2(_04589_),
    .ZN(_05274_));
 AOI221_X2 _22276_ (.A(_05267_),
    .B1(_05269_),
    .B2(net38),
    .C1(_04596_),
    .C2(_05274_),
    .ZN(_05275_));
 INV_X1 _22277_ (.A(_11486_),
    .ZN(_05276_));
 MUX2_X1 _22278_ (.A(_11476_),
    .B(_05276_),
    .S(_11500_),
    .Z(_05277_));
 NOR2_X1 _22279_ (.A1(_04271_),
    .A2(_11505_),
    .ZN(_05278_));
 OAI22_X1 _22280_ (.A1(_04264_),
    .A2(_05277_),
    .B1(_04376_),
    .B2(_05278_),
    .ZN(_05279_));
 AND2_X1 _22281_ (.A1(_11862_),
    .A2(_05279_),
    .ZN(_05280_));
 NOR2_X1 _22282_ (.A1(_15494_),
    .A2(net272),
    .ZN(_05281_));
 NAND4_X2 _22283_ (.A1(_03398_),
    .A2(_03399_),
    .A3(_03415_),
    .A4(_05281_),
    .ZN(_05282_));
 INV_X1 _22284_ (.A(_05241_),
    .ZN(_05283_));
 OR3_X1 _22285_ (.A1(_11482_),
    .A2(_11918_),
    .A3(_05278_),
    .ZN(_05284_));
 OAI33_X1 _22286_ (.A1(_04300_),
    .A2(_11512_),
    .A3(_05278_),
    .B1(_05284_),
    .B2(_04266_),
    .B3(_11510_),
    .ZN(_05285_));
 NOR2_X4 _22287_ (.A1(_04375_),
    .A2(_05285_),
    .ZN(_05286_));
 NAND3_X1 _22288_ (.A1(_05283_),
    .A2(net272),
    .A3(_05286_),
    .ZN(_05287_));
 OAI22_X2 _22289_ (.A1(_05280_),
    .A2(_05282_),
    .B1(_05287_),
    .B2(_03416_),
    .ZN(_05288_));
 AND2_X1 _22290_ (.A1(_03398_),
    .A2(_03399_),
    .ZN(_05289_));
 INV_X1 _22291_ (.A(_15489_),
    .ZN(_05290_));
 AOI21_X2 _22292_ (.A(_03391_),
    .B1(_03219_),
    .B2(_13266_),
    .ZN(_05291_));
 OAI21_X4 _22293_ (.A(_05290_),
    .B1(_05291_),
    .B2(_03418_),
    .ZN(_05292_));
 AND3_X1 _22294_ (.A1(_04264_),
    .A2(_11862_),
    .A3(_04379_),
    .ZN(_05293_));
 NOR3_X1 _22295_ (.A1(_05276_),
    .A2(_04264_),
    .A3(_11918_),
    .ZN(_05294_));
 OAI21_X1 _22296_ (.A(_04273_),
    .B1(_05293_),
    .B2(_05294_),
    .ZN(_05295_));
 NAND3_X1 _22297_ (.A1(_15365_),
    .A2(_04300_),
    .A3(_11862_),
    .ZN(_05296_));
 OAI21_X1 _22298_ (.A(_05295_),
    .B1(_05296_),
    .B2(_04273_),
    .ZN(_05297_));
 OR3_X1 _22299_ (.A1(_05241_),
    .A2(_05292_),
    .A3(_05297_),
    .ZN(_05298_));
 NAND3_X1 _22300_ (.A1(_05283_),
    .A2(_05292_),
    .A3(_05286_),
    .ZN(_05299_));
 AOI21_X1 _22301_ (.A(_05289_),
    .B1(_05298_),
    .B2(_05299_),
    .ZN(_05300_));
 NOR4_X1 _22302_ (.A1(_03412_),
    .A2(_11406_),
    .A3(_03405_),
    .A4(_03411_),
    .ZN(_05301_));
 NOR2_X1 _22303_ (.A1(_11406_),
    .A2(_03413_),
    .ZN(_05302_));
 AOI21_X1 _22304_ (.A(_05301_),
    .B1(_05302_),
    .B2(_03411_),
    .ZN(_05303_));
 OR2_X1 _22305_ (.A1(_04375_),
    .A2(_05285_),
    .ZN(_05304_));
 MUX2_X1 _22306_ (.A(_05304_),
    .B(_05297_),
    .S(net272),
    .Z(_05305_));
 OR3_X1 _22307_ (.A1(_05241_),
    .A2(_05303_),
    .A3(_05305_),
    .ZN(_05306_));
 NOR3_X1 _22308_ (.A1(_11476_),
    .A2(_11918_),
    .A3(_11500_),
    .ZN(_05307_));
 XNOR2_X1 _22309_ (.A(_11482_),
    .B(_11508_),
    .ZN(_05308_));
 OAI22_X1 _22310_ (.A1(_04300_),
    .A2(_11512_),
    .B1(_11918_),
    .B2(_05308_),
    .ZN(_05309_));
 AOI21_X2 _22311_ (.A(_05307_),
    .B1(_05309_),
    .B2(_11505_),
    .ZN(_05310_));
 XNOR2_X2 _22312_ (.A(_15492_),
    .B(_05310_),
    .ZN(_05311_));
 MUX2_X1 _22313_ (.A(_05280_),
    .B(_05304_),
    .S(_05311_),
    .Z(_05312_));
 OAI21_X1 _22314_ (.A(_05306_),
    .B1(_05312_),
    .B2(_05283_),
    .ZN(_05313_));
 OR3_X4 _22315_ (.A1(_05288_),
    .A2(_05300_),
    .A3(_05313_),
    .ZN(_05314_));
 NOR3_X2 _22316_ (.A1(_11918_),
    .A2(_04273_),
    .A3(_04304_),
    .ZN(_05315_));
 INV_X2 _22317_ (.A(_05315_),
    .ZN(_05316_));
 MUX2_X1 _22318_ (.A(_05304_),
    .B(_05280_),
    .S(_05311_),
    .Z(_05317_));
 AND4_X1 _22319_ (.A1(_03398_),
    .A2(_03399_),
    .A3(_03415_),
    .A4(_05281_),
    .ZN(_05318_));
 AOI221_X2 _22320_ (.A(_05315_),
    .B1(_05317_),
    .B2(_15494_),
    .C1(_05304_),
    .C2(_05318_),
    .ZN(_05319_));
 NOR2_X1 _22321_ (.A1(_05241_),
    .A2(_05292_),
    .ZN(_05320_));
 NOR2_X1 _22322_ (.A1(_03415_),
    .A2(_05286_),
    .ZN(_05321_));
 AND4_X1 _22323_ (.A1(_03398_),
    .A2(_03399_),
    .A3(_03415_),
    .A4(_05280_),
    .ZN(_05322_));
 OAI21_X2 _22324_ (.A(_05320_),
    .B1(_05321_),
    .B2(_05322_),
    .ZN(_05323_));
 AOI21_X2 _22325_ (.A(_05286_),
    .B1(_03399_),
    .B2(_03398_),
    .ZN(_05324_));
 AND2_X1 _22326_ (.A1(_05292_),
    .A2(_05280_),
    .ZN(_05325_));
 AOI22_X4 _22327_ (.A1(net273),
    .A2(_05324_),
    .B1(_05325_),
    .B2(_03416_),
    .ZN(_05326_));
 OAI211_X4 _22328_ (.A(_05319_),
    .B(_05323_),
    .C1(_05326_),
    .C2(_05241_),
    .ZN(_05327_));
 INV_X1 _22329_ (.A(\alu_adder_result_ex[10] ),
    .ZN(_05328_));
 NOR4_X1 _22330_ (.A1(\alu_adder_result_ex[16] ),
    .A2(net370),
    .A3(\alu_adder_result_ex[2] ),
    .A4(\alu_adder_result_ex[4] ),
    .ZN(_05329_));
 NAND3_X1 _22331_ (.A1(_05328_),
    .A2(_03417_),
    .A3(_05329_),
    .ZN(_05330_));
 OR4_X2 _22332_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_12949_),
    .A3(_13121_),
    .A4(net382),
    .ZN(_05331_));
 OR3_X1 _22333_ (.A1(\alu_adder_result_ex[13] ),
    .A2(\alu_adder_result_ex[17] ),
    .A3(\alu_adder_result_ex[19] ),
    .ZN(_05332_));
 OR4_X1 _22334_ (.A1(net413),
    .A2(net375),
    .A3(_03623_),
    .A4(_05332_),
    .ZN(_05333_));
 OR4_X1 _22335_ (.A1(\alu_adder_result_ex[15] ),
    .A2(\alu_adder_result_ex[21] ),
    .A3(\alu_adder_result_ex[25] ),
    .A4(net14),
    .ZN(_05334_));
 OR4_X1 _22336_ (.A1(\alu_adder_result_ex[6] ),
    .A2(\alu_adder_result_ex[8] ),
    .A3(_05333_),
    .A4(_05334_),
    .ZN(_05335_));
 OR4_X1 _22337_ (.A1(\alu_adder_result_ex[12] ),
    .A2(\alu_adder_result_ex[14] ),
    .A3(\alu_adder_result_ex[28] ),
    .A4(_05335_),
    .ZN(_05336_));
 NOR4_X2 _22338_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_05330_),
    .A3(_05331_),
    .A4(_05336_),
    .ZN(_05337_));
 MUX2_X2 _22339_ (.A(_05316_),
    .B(_05327_),
    .S(_05337_),
    .Z(_05338_));
 AOI21_X2 _22340_ (.A(_04381_),
    .B1(_05314_),
    .B2(_05338_),
    .ZN(_05339_));
 INV_X1 _22341_ (.A(_15839_),
    .ZN(_05340_));
 AOI22_X1 _22342_ (.A1(_05340_),
    .A2(_04353_),
    .B1(_04368_),
    .B2(\alu_adder_result_ex[0] ),
    .ZN(_05341_));
 AOI22_X1 _22343_ (.A1(_15840_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_15843_),
    .ZN(_05342_));
 OAI21_X1 _22344_ (.A(_05341_),
    .B1(_05342_),
    .B2(_04370_),
    .ZN(_05343_));
 AOI21_X1 _22345_ (.A(_05343_),
    .B1(_05240_),
    .B2(_04840_),
    .ZN(_05344_));
 OAI21_X1 _22346_ (.A(_05344_),
    .B1(_05256_),
    .B2(_04688_),
    .ZN(_05345_));
 OAI221_X2 _22347_ (.A(_04815_),
    .B1(_05339_),
    .B2(_05345_),
    .C1(_10678_),
    .C2(_03465_),
    .ZN(_05346_));
 NOR2_X1 _22348_ (.A1(_15553_),
    .A2(_04625_),
    .ZN(_05347_));
 AOI21_X1 _22349_ (.A(_05347_),
    .B1(_04626_),
    .B2(_00217_),
    .ZN(_05348_));
 NOR2_X2 _22350_ (.A1(_04622_),
    .A2(_05348_),
    .ZN(_05349_));
 NOR2_X1 _22351_ (.A1(_12103_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .ZN(_05350_));
 NOR3_X4 _22352_ (.A1(_11408_),
    .A2(_05349_),
    .A3(_05350_),
    .ZN(_05351_));
 BUF_X2 _22353_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .Z(_05352_));
 AOI22_X2 _22354_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_05352_),
    .ZN(_05353_));
 NOR2_X1 _22355_ (.A1(_04557_),
    .A2(_05353_),
    .ZN(_05354_));
 INV_X1 _22356_ (.A(_00551_),
    .ZN(_05355_));
 INV_X1 _22357_ (.A(_00552_),
    .ZN(_05356_));
 AOI22_X2 _22358_ (.A1(_05355_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_05356_),
    .ZN(_05357_));
 NOR2_X1 _22359_ (.A1(_04559_),
    .A2(_05357_),
    .ZN(_05358_));
 AOI22_X1 _22360_ (.A1(\cs_registers_i.csr_mepc_o[0] ),
    .A2(_05074_),
    .B1(_05228_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .ZN(_05359_));
 AOI22_X1 _22361_ (.A1(\cs_registers_i.mscratch_q[0] ),
    .A2(_04972_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[0] ),
    .ZN(_05360_));
 NAND2_X1 _22362_ (.A1(_05359_),
    .A2(_05360_),
    .ZN(_05361_));
 INV_X1 _22363_ (.A(_00553_),
    .ZN(_05362_));
 AOI22_X1 _22364_ (.A1(_05362_),
    .A2(_05231_),
    .B1(_05198_),
    .B2(\cs_registers_i.dcsr_q[0] ),
    .ZN(_05363_));
 NOR2_X1 _22365_ (.A1(_03530_),
    .A2(_03596_),
    .ZN(_05364_));
 NOR3_X1 _22366_ (.A1(_04251_),
    .A2(_04548_),
    .A3(_05364_),
    .ZN(_05365_));
 AOI221_X1 _22367_ (.A(_05365_),
    .B1(_04526_),
    .B2(net71),
    .C1(\cs_registers_i.dscratch1_q[0] ),
    .C2(_04529_),
    .ZN(_05366_));
 AOI21_X1 _22368_ (.A(_05199_),
    .B1(_04771_),
    .B2(\cs_registers_i.dscratch0_q[0] ),
    .ZN(_05367_));
 NAND3_X1 _22369_ (.A1(_05363_),
    .A2(_05366_),
    .A3(_05367_),
    .ZN(_05368_));
 OR4_X4 _22370_ (.A1(_05354_),
    .A2(_05358_),
    .A3(_05361_),
    .A4(_05368_),
    .ZN(_05369_));
 NOR3_X4 _22371_ (.A1(_04905_),
    .A2(_05351_),
    .A3(_05369_),
    .ZN(_05370_));
 AOI22_X4 _22372_ (.A1(_04611_),
    .A2(_05275_),
    .B1(_05346_),
    .B2(_05370_),
    .ZN(_05371_));
 BUF_X2 _22373_ (.A(_05371_),
    .Z(_05372_));
 NAND2_X2 _22374_ (.A1(_10394_),
    .A2(_11315_),
    .ZN(_05373_));
 NOR2_X4 _22375_ (.A1(_04603_),
    .A2(_05373_),
    .ZN(_05374_));
 NAND2_X4 _22376_ (.A1(_04613_),
    .A2(_05374_),
    .ZN(_05375_));
 BUF_X4 _22377_ (.A(_05375_),
    .Z(_05376_));
 MUX2_X1 _22378_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S(_05376_),
    .Z(_01196_));
 NAND3_X1 _22379_ (.A1(_05268_),
    .A2(_05261_),
    .A3(net46),
    .ZN(_05377_));
 NAND2_X1 _22380_ (.A1(_04594_),
    .A2(net68),
    .ZN(_05378_));
 OAI21_X1 _22381_ (.A(_05377_),
    .B1(_05378_),
    .B2(_04596_),
    .ZN(_05379_));
 NAND2_X1 _22382_ (.A1(_04859_),
    .A2(_05379_),
    .ZN(_05380_));
 AOI22_X1 _22383_ (.A1(\load_store_unit_i.rdata_q[9] ),
    .A2(_05262_),
    .B1(_05265_),
    .B2(\load_store_unit_i.rdata_q[17] ),
    .ZN(_05381_));
 OAI21_X1 _22384_ (.A(_05380_),
    .B1(_05381_),
    .B2(_04859_),
    .ZN(_05382_));
 NAND2_X1 _22385_ (.A1(_05261_),
    .A2(net49),
    .ZN(_05383_));
 NAND2_X2 _22386_ (.A1(_05268_),
    .A2(_04594_),
    .ZN(_05384_));
 AOI22_X2 _22387_ (.A1(_05270_),
    .A2(net54),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[25] ),
    .ZN(_05385_));
 OAI22_X2 _22388_ (.A1(_04597_),
    .A2(_05383_),
    .B1(_05384_),
    .B2(_05385_),
    .ZN(_05386_));
 OAI21_X2 _22389_ (.A(_04611_),
    .B1(_05382_),
    .B2(_05386_),
    .ZN(_05387_));
 NOR2_X1 _22390_ (.A1(_15556_),
    .A2(_04624_),
    .ZN(_05388_));
 AOI21_X2 _22391_ (.A(_05388_),
    .B1(_04624_),
    .B2(_00185_),
    .ZN(_05389_));
 NOR2_X1 _22392_ (.A1(_10310_),
    .A2(_05389_),
    .ZN(_05390_));
 OAI21_X1 _22393_ (.A(_11401_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .B2(_11432_),
    .ZN(_05391_));
 OAI21_X2 _22394_ (.A(_10744_),
    .B1(_05390_),
    .B2(_05391_),
    .ZN(_05392_));
 NAND2_X1 _22395_ (.A1(_15850_),
    .A2(_04353_),
    .ZN(_05393_));
 AOI221_X1 _22396_ (.A(_04351_),
    .B1(_04359_),
    .B2(_15848_),
    .C1(_04983_),
    .C2(_15847_),
    .ZN(_05394_));
 INV_X1 _22397_ (.A(_05394_),
    .ZN(_05395_));
 AOI221_X2 _22398_ (.A(_05392_),
    .B1(_05393_),
    .B2(_05395_),
    .C1(_04369_),
    .C2(net15),
    .ZN(_05396_));
 OAI21_X1 _22399_ (.A(_05396_),
    .B1(_05153_),
    .B2(_04725_),
    .ZN(_05397_));
 NOR2_X1 _22400_ (.A1(_04688_),
    .A2(_05186_),
    .ZN(_05398_));
 NOR2_X1 _22401_ (.A1(_00554_),
    .A2(_04539_),
    .ZN(_05399_));
 AOI221_X2 _22402_ (.A(_05399_),
    .B1(net16),
    .B2(\cs_registers_i.dscratch0_q[1] ),
    .C1(\cs_registers_i.dscratch1_q[1] ),
    .C2(_04775_),
    .ZN(_05400_));
 AOI222_X2 _22403_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(_05022_),
    .B1(_05074_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .C1(\cs_registers_i.mscratch_q[1] ),
    .C2(_04972_),
    .ZN(_05401_));
 AOI222_X2 _22404_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(net17),
    .B1(_05228_),
    .B2(\cs_registers_i.mcause_q[1] ),
    .C1(net82),
    .C2(_04527_),
    .ZN(_05402_));
 AND3_X1 _22405_ (.A1(_05400_),
    .A2(_05401_),
    .A3(_05402_),
    .ZN(_05403_));
 CLKBUF_X3 _22406_ (.A(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .Z(_05404_));
 AOI22_X2 _22407_ (.A1(_05404_),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][33] ),
    .ZN(_05405_));
 AOI22_X2 _22408_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][1] ),
    .ZN(_05406_));
 OAI221_X2 _22409_ (.A(_05403_),
    .B1(_05405_),
    .B2(_05031_),
    .C1(_04560_),
    .C2(_05406_),
    .ZN(_05407_));
 OAI222_X2 _22410_ (.A1(_04815_),
    .A2(_05392_),
    .B1(_05397_),
    .B2(_05398_),
    .C1(_05407_),
    .C2(_04393_),
    .ZN(_05408_));
 OAI21_X2 _22411_ (.A(_05387_),
    .B1(_05408_),
    .B2(_04906_),
    .ZN(_05409_));
 BUF_X2 _22412_ (.A(_05409_),
    .Z(_05410_));
 MUX2_X1 _22413_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .S(_05376_),
    .Z(_01197_));
 BUF_X4 _22414_ (.A(_05093_),
    .Z(_05411_));
 BUF_X4 _22415_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Z(_05412_));
 AOI211_X2 _22416_ (.A(_10899_),
    .B(_05412_),
    .C1(_04605_),
    .C2(_04611_),
    .ZN(_05413_));
 AND2_X1 _22417_ (.A1(_04852_),
    .A2(_05413_),
    .ZN(_05414_));
 BUF_X4 _22418_ (.A(_05414_),
    .Z(_05415_));
 MUX2_X1 _22419_ (.A(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .B(_05411_),
    .S(_05415_),
    .Z(_01198_));
 BUF_X4 _22420_ (.A(_05375_),
    .Z(_05416_));
 NAND2_X1 _22421_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .A2(_05416_),
    .ZN(_05417_));
 AOI22_X1 _22422_ (.A1(_05270_),
    .A2(net55),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[26] ),
    .ZN(_05418_));
 NAND2_X1 _22423_ (.A1(_05261_),
    .A2(net59),
    .ZN(_05419_));
 OAI22_X1 _22424_ (.A1(_05384_),
    .A2(_05418_),
    .B1(_05419_),
    .B2(_04597_),
    .ZN(_05420_));
 CLKBUF_X3 _22425_ (.A(_05268_),
    .Z(_05421_));
 NAND3_X1 _22426_ (.A1(_05421_),
    .A2(_05261_),
    .A3(net47),
    .ZN(_05422_));
 NAND2_X1 _22427_ (.A1(_04594_),
    .A2(net39),
    .ZN(_05423_));
 OAI221_X1 _22428_ (.A(_05422_),
    .B1(_05423_),
    .B2(_05421_),
    .C1(_04574_),
    .C2(_05270_),
    .ZN(_05424_));
 AOI22_X1 _22429_ (.A1(\load_store_unit_i.rdata_q[10] ),
    .A2(_05262_),
    .B1(_05265_),
    .B2(\load_store_unit_i.rdata_q[18] ),
    .ZN(_05425_));
 NAND2_X1 _22430_ (.A1(_04582_),
    .A2(_05425_),
    .ZN(_05426_));
 AOI21_X1 _22431_ (.A(_05420_),
    .B1(_05424_),
    .B2(_05426_),
    .ZN(_05427_));
 OR2_X1 _22432_ (.A1(_00556_),
    .A2(_04463_),
    .ZN(_05428_));
 NAND2_X1 _22433_ (.A1(_15565_),
    .A2(_04463_),
    .ZN(_05429_));
 NAND3_X2 _22434_ (.A1(_12102_),
    .A2(_05428_),
    .A3(_05429_),
    .ZN(_05430_));
 INV_X1 _22435_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .ZN(_05431_));
 AOI21_X2 _22436_ (.A(_11407_),
    .B1(_05431_),
    .B2(net304),
    .ZN(_05432_));
 AOI22_X1 _22437_ (.A1(_15855_),
    .A2(_04360_),
    .B1(_04983_),
    .B2(_15854_),
    .ZN(_05433_));
 MUX2_X1 _22438_ (.A(_15858_),
    .B(_05433_),
    .S(_04664_),
    .Z(_05434_));
 NAND2_X1 _22439_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_04368_),
    .ZN(_05435_));
 NAND2_X1 _22440_ (.A1(_05434_),
    .A2(_05435_),
    .ZN(_05436_));
 AOI221_X2 _22441_ (.A(_04662_),
    .B1(_05430_),
    .B2(_05432_),
    .C1(_05436_),
    .C2(_04815_),
    .ZN(_05437_));
 NOR2_X1 _22442_ (.A1(_04987_),
    .A2(_05007_),
    .ZN(_05438_));
 NAND2_X1 _22443_ (.A1(_04840_),
    .A2(_04816_),
    .ZN(_05439_));
 NAND3_X1 _22444_ (.A1(_05128_),
    .A2(_05131_),
    .A3(_05132_),
    .ZN(_05440_));
 OAI221_X2 _22445_ (.A(_05437_),
    .B1(_05438_),
    .B2(_05439_),
    .C1(_05440_),
    .C2(_04688_),
    .ZN(_05441_));
 AOI22_X1 _22446_ (.A1(\cs_registers_i.mtval_q[2] ),
    .A2(_05022_),
    .B1(_05228_),
    .B2(\cs_registers_i.mcause_q[2] ),
    .ZN(_05442_));
 AOI22_X1 _22447_ (.A1(\cs_registers_i.mscratch_q[2] ),
    .A2(_04972_),
    .B1(_05074_),
    .B2(\cs_registers_i.csr_mepc_o[2] ),
    .ZN(_05443_));
 NAND2_X1 _22448_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_04773_),
    .ZN(_05444_));
 OR3_X1 _22449_ (.A1(_03496_),
    .A2(_04251_),
    .A3(_04730_),
    .ZN(_05445_));
 INV_X1 _22450_ (.A(_01162_),
    .ZN(_05446_));
 AOI22_X1 _22451_ (.A1(\cs_registers_i.dscratch0_q[2] ),
    .A2(_04510_),
    .B1(_05198_),
    .B2(_05446_),
    .ZN(_05447_));
 AND3_X1 _22452_ (.A1(_05444_),
    .A2(_05445_),
    .A3(_05447_),
    .ZN(_05448_));
 INV_X1 _22453_ (.A(\cs_registers_i.dscratch1_q[2] ),
    .ZN(_05449_));
 OAI211_X2 _22454_ (.A(_03506_),
    .B(_04538_),
    .C1(_03530_),
    .C2(_10920_),
    .ZN(_05450_));
 OAI21_X1 _22455_ (.A(_10922_),
    .B1(_03513_),
    .B2(_03524_),
    .ZN(_05451_));
 NAND2_X2 _22456_ (.A1(_04239_),
    .A2(_05451_),
    .ZN(_05452_));
 OAI22_X1 _22457_ (.A1(_05449_),
    .A2(_05450_),
    .B1(_05452_),
    .B2(_04735_),
    .ZN(_05453_));
 INV_X1 _22458_ (.A(_01159_),
    .ZN(_05454_));
 AOI221_X1 _22459_ (.A(_05453_),
    .B1(_04527_),
    .B2(net93),
    .C1(_05454_),
    .C2(_05231_),
    .ZN(_05455_));
 AND4_X1 _22460_ (.A1(_05442_),
    .A2(_05443_),
    .A3(_05448_),
    .A4(_05455_),
    .ZN(_05456_));
 CLKBUF_X3 _22461_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .Z(_05457_));
 AOI22_X2 _22462_ (.A1(_05457_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][34] ),
    .ZN(_05458_));
 BUF_X2 _22463_ (.A(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .Z(_05459_));
 AOI22_X2 _22464_ (.A1(_05459_),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][2] ),
    .ZN(_05460_));
 OAI221_X2 _22465_ (.A(_05456_),
    .B1(_05458_),
    .B2(_04557_),
    .C1(_04783_),
    .C2(_05460_),
    .ZN(_05461_));
 OAI21_X2 _22466_ (.A(_05441_),
    .B1(_05461_),
    .B2(_04563_),
    .ZN(_05462_));
 MUX2_X1 _22467_ (.A(_05427_),
    .B(_05462_),
    .S(_04600_),
    .Z(_05463_));
 CLKBUF_X3 _22468_ (.A(_05463_),
    .Z(_05464_));
 BUF_X4 _22469_ (.A(_05375_),
    .Z(_05465_));
 OAI21_X1 _22470_ (.A(_05417_),
    .B1(_05464_),
    .B2(_05465_),
    .ZN(_01199_));
 NAND2_X1 _22471_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .A2(_05416_),
    .ZN(_05466_));
 NOR2_X1 _22472_ (.A1(_15580_),
    .A2(_04624_),
    .ZN(_05467_));
 AOI21_X1 _22473_ (.A(_05467_),
    .B1(_04625_),
    .B2(_00557_),
    .ZN(_05468_));
 NOR2_X2 _22474_ (.A1(_10310_),
    .A2(_05468_),
    .ZN(_05469_));
 OAI21_X1 _22475_ (.A(_11401_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .B2(_11432_),
    .ZN(_05470_));
 AOI221_X1 _22476_ (.A(_04350_),
    .B1(_04358_),
    .B2(_15863_),
    .C1(_04361_),
    .C2(_15866_),
    .ZN(_05471_));
 AOI21_X1 _22477_ (.A(_05471_),
    .B1(_04352_),
    .B2(_15862_),
    .ZN(_05472_));
 AOI21_X1 _22478_ (.A(_05472_),
    .B1(_04368_),
    .B2(\alu_adder_result_ex[3] ),
    .ZN(_05473_));
 OAI22_X1 _22479_ (.A1(_05469_),
    .A2(_05470_),
    .B1(_05473_),
    .B2(_04389_),
    .ZN(_05474_));
 AND3_X2 _22480_ (.A1(_04279_),
    .A2(_04280_),
    .A3(_04306_),
    .ZN(_05475_));
 NAND2_X1 _22481_ (.A1(_04456_),
    .A2(_05475_),
    .ZN(_05476_));
 NAND2_X1 _22482_ (.A1(_04393_),
    .A2(_05476_),
    .ZN(_05477_));
 OR2_X1 _22483_ (.A1(_05474_),
    .A2(_05477_),
    .ZN(_05478_));
 AOI21_X1 _22484_ (.A(_04458_),
    .B1(_04830_),
    .B2(_04720_),
    .ZN(_05479_));
 NOR2_X2 _22485_ (.A1(_04342_),
    .A2(_04281_),
    .ZN(_05480_));
 AOI221_X2 _22486_ (.A(_05478_),
    .B1(_05479_),
    .B2(_05480_),
    .C1(_05056_),
    .C2(_04276_),
    .ZN(_05481_));
 CLKBUF_X3 _22487_ (.A(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .Z(_05482_));
 BUF_X2 _22488_ (.A(\cs_registers_i.mhpmcounter[2][35] ),
    .Z(_05483_));
 AOI22_X2 _22489_ (.A1(_05482_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_05483_),
    .ZN(_05484_));
 NOR2_X1 _22490_ (.A1(_04557_),
    .A2(_05484_),
    .ZN(_05485_));
 AOI22_X1 _22491_ (.A1(\cs_registers_i.csr_mepc_o[3] ),
    .A2(_05074_),
    .B1(_05228_),
    .B2(\cs_registers_i.mcause_q[3] ),
    .ZN(_05486_));
 NOR2_X4 _22492_ (.A1(_11072_),
    .A2(_05452_),
    .ZN(_05487_));
 AOI222_X2 _22493_ (.A1(\cs_registers_i.dscratch0_q[3] ),
    .A2(net16),
    .B1(_04529_),
    .B2(\cs_registers_i.dscratch1_q[3] ),
    .C1(\cs_registers_i.csr_mstatus_mie_o ),
    .C2(_05487_),
    .ZN(_05488_));
 NAND4_X2 _22494_ (.A1(_15869_),
    .A2(_03491_),
    .A3(_03485_),
    .A4(_03514_),
    .ZN(_05489_));
 NOR2_X2 _22495_ (.A1(_03575_),
    .A2(_05489_),
    .ZN(_05490_));
 AOI222_X2 _22496_ (.A1(\cs_registers_i.mie_q[17] ),
    .A2(_04514_),
    .B1(_04773_),
    .B2(_03950_),
    .C1(net96),
    .C2(_05490_),
    .ZN(_05491_));
 NAND4_X1 _22497_ (.A1(_04534_),
    .A2(_05486_),
    .A3(_05488_),
    .A4(_05491_),
    .ZN(_05492_));
 AOI222_X2 _22498_ (.A1(net151),
    .A2(_04517_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[3] ),
    .C1(\cs_registers_i.mscratch_q[3] ),
    .C2(_04523_),
    .ZN(_05493_));
 BUF_X2 _22499_ (.A(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .Z(_05494_));
 AOI22_X2 _22500_ (.A1(_05494_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\cs_registers_i.mhpmcounter[2][3] ),
    .ZN(_05495_));
 OAI21_X1 _22501_ (.A(_05493_),
    .B1(_05495_),
    .B2(_04559_),
    .ZN(_05496_));
 OR3_X2 _22502_ (.A1(_05485_),
    .A2(_05492_),
    .A3(_05496_),
    .ZN(_05497_));
 NOR2_X1 _22503_ (.A1(_04563_),
    .A2(_05497_),
    .ZN(_05498_));
 OAI21_X1 _22504_ (.A(_04764_),
    .B1(_05481_),
    .B2(_05498_),
    .ZN(_05499_));
 AOI22_X1 _22505_ (.A1(\load_store_unit_i.rdata_q[11] ),
    .A2(_05262_),
    .B1(_05265_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .ZN(_05500_));
 NOR2_X1 _22506_ (.A1(_04859_),
    .A2(_05500_),
    .ZN(_05501_));
 NAND3_X1 _22507_ (.A1(_04596_),
    .A2(_05261_),
    .A3(net48),
    .ZN(_05502_));
 NAND2_X1 _22508_ (.A1(_04594_),
    .A2(net40),
    .ZN(_05503_));
 OAI21_X1 _22509_ (.A(_05502_),
    .B1(_05503_),
    .B2(_04596_),
    .ZN(_05504_));
 AOI21_X1 _22510_ (.A(_05501_),
    .B1(_05504_),
    .B2(_04859_),
    .ZN(_05505_));
 AOI22_X2 _22511_ (.A1(_05270_),
    .A2(net56),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[27] ),
    .ZN(_05506_));
 NAND2_X1 _22512_ (.A1(_05261_),
    .A2(net62),
    .ZN(_05507_));
 OAI221_X2 _22513_ (.A(_05505_),
    .B1(_05506_),
    .B2(_05384_),
    .C1(_05507_),
    .C2(_04597_),
    .ZN(_05508_));
 OAI21_X2 _22514_ (.A(_05499_),
    .B1(_05508_),
    .B2(_04764_),
    .ZN(_05509_));
 CLKBUF_X3 _22515_ (.A(_05509_),
    .Z(_05510_));
 OAI21_X1 _22516_ (.A(_05466_),
    .B1(_05510_),
    .B2(_05465_),
    .ZN(_01200_));
 AOI22_X1 _22517_ (.A1(\load_store_unit_i.rdata_q[12] ),
    .A2(_05262_),
    .B1(_05265_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .ZN(_05511_));
 NOR2_X1 _22518_ (.A1(_04859_),
    .A2(_05511_),
    .ZN(_05512_));
 CLKBUF_X3 _22519_ (.A(_04570_),
    .Z(_05513_));
 NAND3_X1 _22520_ (.A1(_05513_),
    .A2(_04589_),
    .A3(net50),
    .ZN(_05514_));
 NAND2_X1 _22521_ (.A1(_04586_),
    .A2(net41),
    .ZN(_05515_));
 OAI21_X1 _22522_ (.A(_05514_),
    .B1(_05515_),
    .B2(_05268_),
    .ZN(_05516_));
 AOI21_X1 _22523_ (.A(_05512_),
    .B1(_05516_),
    .B2(_04859_),
    .ZN(_05517_));
 AOI22_X2 _22524_ (.A1(_05270_),
    .A2(net57),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[28] ),
    .ZN(_05518_));
 NAND2_X1 _22525_ (.A1(_05261_),
    .A2(net63),
    .ZN(_05519_));
 OAI221_X2 _22526_ (.A(_05517_),
    .B1(_05518_),
    .B2(_05384_),
    .C1(_05519_),
    .C2(_04597_),
    .ZN(_05520_));
 NOR2_X1 _22527_ (.A1(_15588_),
    .A2(_04624_),
    .ZN(_05521_));
 AOI21_X1 _22528_ (.A(_05521_),
    .B1(_04624_),
    .B2(_00558_),
    .ZN(_05522_));
 NOR2_X2 _22529_ (.A1(_10310_),
    .A2(_05522_),
    .ZN(_05523_));
 OAI21_X1 _22530_ (.A(_11401_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B2(_11432_),
    .ZN(_05524_));
 AOI221_X2 _22531_ (.A(_04350_),
    .B1(_04358_),
    .B2(_15871_),
    .C1(_04361_),
    .C2(_15870_),
    .ZN(_05525_));
 AOI21_X1 _22532_ (.A(_05525_),
    .B1(_04352_),
    .B2(_15874_),
    .ZN(_05526_));
 AOI21_X1 _22533_ (.A(_05526_),
    .B1(_04368_),
    .B2(\alu_adder_result_ex[4] ),
    .ZN(_05527_));
 OAI221_X2 _22534_ (.A(_10744_),
    .B1(_05523_),
    .B2(_05524_),
    .C1(_05527_),
    .C2(_04390_),
    .ZN(_05528_));
 AND2_X1 _22535_ (.A1(_04840_),
    .A2(_04816_),
    .ZN(_05529_));
 AOI221_X2 _22536_ (.A(_05528_),
    .B1(_05529_),
    .B2(_04821_),
    .C1(_04276_),
    .C2(_04846_),
    .ZN(_05530_));
 AOI222_X2 _22537_ (.A1(\cs_registers_i.mtval_q[4] ),
    .A2(_05022_),
    .B1(_05074_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .C1(_05228_),
    .C2(\cs_registers_i.mcause_q[4] ),
    .ZN(_05531_));
 NOR2_X1 _22538_ (.A1(_01164_),
    .A2(_04539_),
    .ZN(_05532_));
 AOI221_X1 _22539_ (.A(_05532_),
    .B1(_04510_),
    .B2(\cs_registers_i.dscratch0_q[4] ),
    .C1(\cs_registers_i.dscratch1_q[4] ),
    .C2(_04529_),
    .ZN(_05533_));
 AOI221_X1 _22540_ (.A(_05231_),
    .B1(_04527_),
    .B2(net97),
    .C1(\cs_registers_i.mscratch_q[4] ),
    .C2(_04523_),
    .ZN(_05534_));
 AND3_X1 _22541_ (.A1(_05531_),
    .A2(_05533_),
    .A3(_05534_),
    .ZN(_05535_));
 BUF_X2 _22542_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .Z(_05536_));
 AOI22_X2 _22543_ (.A1(_05536_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][36] ),
    .ZN(_05537_));
 BUF_X1 _22544_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .Z(_05538_));
 AOI22_X2 _22545_ (.A1(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(_05538_),
    .ZN(_05539_));
 OAI221_X2 _22546_ (.A(_05535_),
    .B1(_05537_),
    .B2(_05031_),
    .C1(_04783_),
    .C2(_05539_),
    .ZN(_05540_));
 NOR2_X1 _22547_ (.A1(_04393_),
    .A2(_05540_),
    .ZN(_05541_));
 NOR2_X2 _22548_ (.A1(_05530_),
    .A2(_05541_),
    .ZN(_05542_));
 MUX2_X2 _22549_ (.A(_05520_),
    .B(_05542_),
    .S(_04263_),
    .Z(_05543_));
 BUF_X2 _22550_ (.A(_05543_),
    .Z(_05544_));
 MUX2_X1 _22551_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .S(_05376_),
    .Z(_01201_));
 AOI22_X1 _22552_ (.A1(\load_store_unit_i.rdata_q[13] ),
    .A2(_05262_),
    .B1(_05265_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .ZN(_05545_));
 NOR2_X1 _22553_ (.A1(_04858_),
    .A2(_05545_),
    .ZN(_05546_));
 NAND3_X1 _22554_ (.A1(_05513_),
    .A2(_04589_),
    .A3(net51),
    .ZN(_05547_));
 NAND2_X1 _22555_ (.A1(_04586_),
    .A2(net42),
    .ZN(_05548_));
 OAI21_X1 _22556_ (.A(_05547_),
    .B1(_05548_),
    .B2(_05268_),
    .ZN(_05549_));
 AOI21_X1 _22557_ (.A(_05546_),
    .B1(_05549_),
    .B2(_04859_),
    .ZN(_05550_));
 AOI22_X2 _22558_ (.A1(_05270_),
    .A2(net58),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[29] ),
    .ZN(_05551_));
 NAND2_X1 _22559_ (.A1(_05261_),
    .A2(net64),
    .ZN(_05552_));
 OAI221_X2 _22560_ (.A(_05550_),
    .B1(_05551_),
    .B2(_05384_),
    .C1(_05552_),
    .C2(_04597_),
    .ZN(_05553_));
 NOR2_X1 _22561_ (.A1(_14126_),
    .A2(_04625_),
    .ZN(_05554_));
 AOI21_X1 _22562_ (.A(_05554_),
    .B1(_05079_),
    .B2(_00559_),
    .ZN(_05555_));
 NOR2_X2 _22563_ (.A1(_04622_),
    .A2(_05555_),
    .ZN(_05556_));
 OAI21_X1 _22564_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B2(_12102_),
    .ZN(_05557_));
 OAI21_X2 _22565_ (.A(_04393_),
    .B1(_05556_),
    .B2(_05557_),
    .ZN(_05558_));
 MUX2_X1 _22566_ (.A(_15879_),
    .B(_15878_),
    .S(_04983_),
    .Z(_05559_));
 NAND2_X1 _22567_ (.A1(_04665_),
    .A2(_05559_),
    .ZN(_05560_));
 OAI21_X1 _22568_ (.A(_05560_),
    .B1(_04665_),
    .B2(_15882_),
    .ZN(_05561_));
 INV_X2 _22569_ (.A(_04387_),
    .ZN(_05562_));
 AOI22_X1 _22570_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_04825_),
    .B1(_05561_),
    .B2(_05562_),
    .ZN(_05563_));
 NAND2_X1 _22571_ (.A1(_04457_),
    .A2(_04816_),
    .ZN(_05564_));
 OAI21_X1 _22572_ (.A(_05563_),
    .B1(_05564_),
    .B2(_04991_),
    .ZN(_05565_));
 AOI21_X2 _22573_ (.A(_05558_),
    .B1(_05565_),
    .B2(_04815_),
    .ZN(_05566_));
 NAND2_X1 _22574_ (.A1(_04276_),
    .A2(_05019_),
    .ZN(_05567_));
 AOI22_X2 _22575_ (.A1(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][37] ),
    .ZN(_05568_));
 NOR2_X1 _22576_ (.A1(_05031_),
    .A2(_05568_),
    .ZN(_05569_));
 AOI22_X1 _22577_ (.A1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(\cs_registers_i.mhpmcounter[2][5] ),
    .ZN(_05570_));
 NOR2_X1 _22578_ (.A1(_04559_),
    .A2(_05570_),
    .ZN(_05571_));
 AOI22_X1 _22579_ (.A1(\cs_registers_i.mscratch_q[5] ),
    .A2(_04524_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[5] ),
    .ZN(_05572_));
 AOI221_X2 _22580_ (.A(_05231_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .C1(\cs_registers_i.dscratch0_q[5] ),
    .C2(net16),
    .ZN(_05573_));
 NOR2_X1 _22581_ (.A1(_01165_),
    .A2(_04539_),
    .ZN(_05574_));
 AOI221_X2 _22582_ (.A(_05574_),
    .B1(_04527_),
    .B2(net98),
    .C1(\cs_registers_i.dscratch1_q[5] ),
    .C2(_04529_),
    .ZN(_05575_));
 NAND3_X2 _22583_ (.A1(_05572_),
    .A2(_05573_),
    .A3(_05575_),
    .ZN(_05576_));
 NOR3_X4 _22584_ (.A1(_05569_),
    .A2(_05571_),
    .A3(_05576_),
    .ZN(_05577_));
 AOI22_X4 _22585_ (.A1(_05566_),
    .A2(_05567_),
    .B1(_05577_),
    .B2(_04662_),
    .ZN(_05578_));
 MUX2_X2 _22586_ (.A(_05553_),
    .B(_05578_),
    .S(_04263_),
    .Z(_05579_));
 BUF_X2 _22587_ (.A(_05579_),
    .Z(_05580_));
 MUX2_X1 _22588_ (.A(_05580_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .S(_05376_),
    .Z(_01202_));
 AOI221_X1 _22589_ (.A(_04581_),
    .B1(_04592_),
    .B2(_04570_),
    .C1(_05262_),
    .C2(net43),
    .ZN(_05581_));
 AOI221_X1 _22590_ (.A(_04858_),
    .B1(_05262_),
    .B2(\load_store_unit_i.rdata_q[14] ),
    .C1(_05265_),
    .C2(\load_store_unit_i.rdata_q[22] ),
    .ZN(_05582_));
 OR2_X1 _22591_ (.A1(_05581_),
    .A2(_05582_),
    .ZN(_05583_));
 AOI22_X1 _22592_ (.A1(_05270_),
    .A2(net60),
    .B1(_05272_),
    .B2(\load_store_unit_i.rdata_q[30] ),
    .ZN(_05584_));
 OAI21_X1 _22593_ (.A(_05583_),
    .B1(_05584_),
    .B2(_05261_),
    .ZN(_05585_));
 AOI21_X1 _22594_ (.A(_04587_),
    .B1(_05583_),
    .B2(_04594_),
    .ZN(_05586_));
 MUX2_X1 _22595_ (.A(_05585_),
    .B(_05586_),
    .S(_04619_),
    .Z(_05587_));
 NAND2_X1 _22596_ (.A1(_04611_),
    .A2(_05587_),
    .ZN(_05588_));
 NAND2_X1 _22597_ (.A1(_00560_),
    .A2(_05079_),
    .ZN(_05589_));
 NAND2_X1 _22598_ (.A1(_04461_),
    .A2(_04502_),
    .ZN(_05590_));
 AOI21_X2 _22599_ (.A(_10493_),
    .B1(_05589_),
    .B2(_05590_),
    .ZN(_05591_));
 OAI21_X1 _22600_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B2(_12102_),
    .ZN(_05592_));
 AOI221_X2 _22601_ (.A(_04351_),
    .B1(_04359_),
    .B2(_15887_),
    .C1(_04983_),
    .C2(_15886_),
    .ZN(_05593_));
 AOI21_X1 _22602_ (.A(_05593_),
    .B1(_04370_),
    .B2(_15890_),
    .ZN(_05594_));
 AOI21_X1 _22603_ (.A(_05594_),
    .B1(_04825_),
    .B2(\alu_adder_result_ex[6] ),
    .ZN(_05595_));
 OAI221_X1 _22604_ (.A(_04393_),
    .B1(_05591_),
    .B2(_05592_),
    .C1(_05595_),
    .C2(_04390_),
    .ZN(_05596_));
 INV_X1 _22605_ (.A(_05596_),
    .ZN(_05597_));
 OAI221_X2 _22606_ (.A(_05597_),
    .B1(_05439_),
    .B2(_04952_),
    .C1(_04688_),
    .C2(_04939_),
    .ZN(_05598_));
 AOI221_X1 _22607_ (.A(_04741_),
    .B1(_04743_),
    .B2(net99),
    .C1(\cs_registers_i.mtval_q[6] ),
    .C2(_04747_),
    .ZN(_05599_));
 AOI22_X1 _22608_ (.A1(\cs_registers_i.mscratch_q[6] ),
    .A2(_04738_),
    .B1(_04749_),
    .B2(\cs_registers_i.dscratch1_q[6] ),
    .ZN(_05600_));
 INV_X1 _22609_ (.A(_01166_),
    .ZN(_05601_));
 NOR2_X1 _22610_ (.A1(_11072_),
    .A2(_03498_),
    .ZN(_05602_));
 AOI22_X1 _22611_ (.A1(_05601_),
    .A2(_04736_),
    .B1(_05602_),
    .B2(\cs_registers_i.dcsr_q[6] ),
    .ZN(_05603_));
 AOI22_X1 _22612_ (.A1(\cs_registers_i.dscratch0_q[6] ),
    .A2(_04731_),
    .B1(_04748_),
    .B2(\cs_registers_i.csr_mepc_o[6] ),
    .ZN(_05604_));
 AND4_X1 _22613_ (.A1(_05599_),
    .A2(_05600_),
    .A3(_05603_),
    .A4(_05604_),
    .ZN(_05605_));
 CLKBUF_X2 _22614_ (.A(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .Z(_05606_));
 CLKBUF_X2 _22615_ (.A(\cs_registers_i.mhpmcounter[2][6] ),
    .Z(_05607_));
 AOI22_X2 _22616_ (.A1(_05606_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(_05607_),
    .ZN(_05608_));
 BUF_X2 _22617_ (.A(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .Z(_05609_));
 AOI22_X4 _22618_ (.A1(_05609_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][38] ),
    .ZN(_05610_));
 OAI221_X2 _22619_ (.A(_05605_),
    .B1(_05608_),
    .B2(_03532_),
    .C1(_04756_),
    .C2(_05610_),
    .ZN(_05611_));
 OAI21_X2 _22620_ (.A(_05598_),
    .B1(_05611_),
    .B2(_04563_),
    .ZN(_05612_));
 OAI21_X4 _22621_ (.A(_05588_),
    .B1(_05612_),
    .B2(_04906_),
    .ZN(_05613_));
 BUF_X2 _22622_ (.A(_05613_),
    .Z(_05614_));
 MUX2_X1 _22623_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S(_05376_),
    .Z(_01203_));
 NOR2_X1 _22624_ (.A1(_04585_),
    .A2(_04573_),
    .ZN(_05615_));
 AOI22_X1 _22625_ (.A1(_04593_),
    .A2(\load_store_unit_i.rdata_q[31] ),
    .B1(\load_store_unit_i.rdata_q[23] ),
    .B2(_05615_),
    .ZN(_05616_));
 AOI221_X1 _22626_ (.A(_04589_),
    .B1(_04573_),
    .B2(\load_store_unit_i.rdata_q[31] ),
    .C1(net61),
    .C2(_04565_),
    .ZN(_05617_));
 AOI21_X1 _22627_ (.A(_04593_),
    .B1(_04568_),
    .B2(_04858_),
    .ZN(_05618_));
 OAI22_X1 _22628_ (.A1(_05270_),
    .A2(_05616_),
    .B1(_05617_),
    .B2(_05618_),
    .ZN(_05619_));
 MUX2_X1 _22629_ (.A(\load_store_unit_i.rdata_q[15] ),
    .B(net44),
    .S(_04858_),
    .Z(_05620_));
 MUX2_X1 _22630_ (.A(net66),
    .B(_05620_),
    .S(_04593_),
    .Z(_05621_));
 MUX2_X1 _22631_ (.A(_05619_),
    .B(_05621_),
    .S(_04619_),
    .Z(_05622_));
 NOR2_X2 _22632_ (.A1(_04263_),
    .A2(_05622_),
    .ZN(_05623_));
 AOI21_X2 _22633_ (.A(_04688_),
    .B1(_04876_),
    .B2(_04884_),
    .ZN(_05624_));
 CLKBUF_X3 _22634_ (.A(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .Z(_05625_));
 AOI22_X2 _22635_ (.A1(_05625_),
    .A2(_04550_),
    .B1(_04553_),
    .B2(\cs_registers_i.mhpmcounter[2][39] ),
    .ZN(_05626_));
 NOR2_X1 _22636_ (.A1(_04557_),
    .A2(_05626_),
    .ZN(_05627_));
 CLKBUF_X2 _22637_ (.A(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .Z(_05628_));
 AOI22_X2 _22638_ (.A1(_05628_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\cs_registers_i.mhpmcounter[2][7] ),
    .ZN(_05629_));
 NOR2_X1 _22639_ (.A1(_04559_),
    .A2(_05629_),
    .ZN(_05630_));
 AOI22_X1 _22640_ (.A1(net152),
    .A2(_04518_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[7] ),
    .ZN(_05631_));
 AOI22_X1 _22641_ (.A1(\cs_registers_i.mscratch_q[7] ),
    .A2(_04524_),
    .B1(_05074_),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .ZN(_05632_));
 NAND2_X1 _22642_ (.A1(_05631_),
    .A2(_05632_),
    .ZN(_05633_));
 AOI22_X1 _22643_ (.A1(\cs_registers_i.dscratch0_q[7] ),
    .A2(_04771_),
    .B1(net17),
    .B2(\cs_registers_i.dcsr_q[7] ),
    .ZN(_05634_));
 AOI21_X1 _22644_ (.A(_05231_),
    .B1(_04775_),
    .B2(\cs_registers_i.dscratch1_q[7] ),
    .ZN(_05635_));
 NAND2_X1 _22645_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_04773_),
    .ZN(_05636_));
 AOI222_X2 _22646_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(_04514_),
    .B1(_05487_),
    .B2(\cs_registers_i.mstack_d[2] ),
    .C1(net100),
    .C2(_05490_),
    .ZN(_05637_));
 NAND4_X2 _22647_ (.A1(_05634_),
    .A2(_05635_),
    .A3(_05636_),
    .A4(_05637_),
    .ZN(_05638_));
 OR4_X4 _22648_ (.A1(_05627_),
    .A2(_05630_),
    .A3(_05633_),
    .A4(_05638_),
    .ZN(_05639_));
 MUX2_X1 _22649_ (.A(_15895_),
    .B(_15894_),
    .S(_04363_),
    .Z(_05640_));
 NAND2_X1 _22650_ (.A1(_04665_),
    .A2(_05640_),
    .ZN(_05641_));
 OAI21_X1 _22651_ (.A(_05641_),
    .B1(_04665_),
    .B2(_15898_),
    .ZN(_05642_));
 AOI22_X1 _22652_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_04825_),
    .B1(_05642_),
    .B2(_05562_),
    .ZN(_05643_));
 NAND2_X1 _22653_ (.A1(_04867_),
    .A2(_05529_),
    .ZN(_05644_));
 AOI21_X2 _22654_ (.A(_04391_),
    .B1(_05643_),
    .B2(_05644_),
    .ZN(_05645_));
 NOR2_X1 _22655_ (.A1(_05079_),
    .A2(_04631_),
    .ZN(_05646_));
 AOI21_X1 _22656_ (.A(_05646_),
    .B1(_04626_),
    .B2(_00561_),
    .ZN(_05647_));
 NOR2_X1 _22657_ (.A1(net304),
    .A2(_05647_),
    .ZN(_05648_));
 OAI21_X1 _22658_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B2(_12103_),
    .ZN(_05649_));
 NOR2_X2 _22659_ (.A1(_05648_),
    .A2(_05649_),
    .ZN(_05650_));
 NOR4_X4 _22660_ (.A1(_05624_),
    .A2(_05639_),
    .A3(_05645_),
    .A4(_05650_),
    .ZN(_05651_));
 AOI21_X4 _22661_ (.A(_05623_),
    .B1(_05651_),
    .B2(_04600_),
    .ZN(_05652_));
 BUF_X2 _22662_ (.A(_05652_),
    .Z(_05653_));
 MUX2_X1 _22663_ (.A(_05653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .S(_05376_),
    .Z(_01204_));
 NAND2_X1 _22664_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .A2(_05416_),
    .ZN(_05654_));
 MUX2_X1 _22665_ (.A(_04860_),
    .B(_04862_),
    .S(_05268_),
    .Z(_05655_));
 MUX2_X1 _22666_ (.A(net67),
    .B(\load_store_unit_i.rdata_q[16] ),
    .S(_04585_),
    .Z(_05656_));
 MUX2_X1 _22667_ (.A(\load_store_unit_i.rdata_q[24] ),
    .B(net38),
    .S(_04585_),
    .Z(_05657_));
 MUX2_X1 _22668_ (.A(_05656_),
    .B(_05657_),
    .S(_05268_),
    .Z(_05658_));
 AOI22_X2 _22669_ (.A1(_04574_),
    .A2(_05655_),
    .B1(_05658_),
    .B2(_04582_),
    .ZN(_05659_));
 AOI21_X2 _22670_ (.A(_04263_),
    .B1(_04572_),
    .B2(_05659_),
    .ZN(_05660_));
 AOI21_X4 _22671_ (.A(_03493_),
    .B1(_04456_),
    .B2(_05475_),
    .ZN(_05661_));
 NOR2_X1 _22672_ (.A1(_00562_),
    .A2(_04463_),
    .ZN(_05662_));
 NOR2_X1 _22673_ (.A1(_04624_),
    .A2(_04886_),
    .ZN(_05663_));
 NOR3_X4 _22674_ (.A1(_10310_),
    .A2(_05662_),
    .A3(_05663_),
    .ZN(_05664_));
 OAI21_X1 _22675_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B2(_11432_),
    .ZN(_05665_));
 MUX2_X1 _22676_ (.A(_15903_),
    .B(_15902_),
    .S(_04362_),
    .Z(_05666_));
 NAND2_X1 _22677_ (.A1(_04664_),
    .A2(_05666_),
    .ZN(_05667_));
 OAI21_X1 _22678_ (.A(_05667_),
    .B1(_04664_),
    .B2(_15906_),
    .ZN(_05668_));
 AOI22_X2 _22679_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_04368_),
    .B1(_05668_),
    .B2(_05562_),
    .ZN(_05669_));
 OAI221_X2 _22680_ (.A(_05661_),
    .B1(_05664_),
    .B2(_05665_),
    .C1(_05669_),
    .C2(_04390_),
    .ZN(_05670_));
 NOR2_X1 _22681_ (.A1(_04725_),
    .A2(_04987_),
    .ZN(_05671_));
 AOI221_X2 _22682_ (.A(_05670_),
    .B1(_05671_),
    .B2(_04684_),
    .C1(_04457_),
    .C2(_04678_),
    .ZN(_05672_));
 OR2_X1 _22683_ (.A1(_04688_),
    .A2(_04724_),
    .ZN(_05673_));
 AOI222_X2 _22684_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(_04521_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[8] ),
    .C1(\cs_registers_i.mscratch_q[8] ),
    .C2(_04524_),
    .ZN(_05674_));
 INV_X1 _22685_ (.A(_05674_),
    .ZN(_05675_));
 AOI22_X2 _22686_ (.A1(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][40] ),
    .ZN(_05676_));
 NOR2_X2 _22687_ (.A1(_05031_),
    .A2(_05676_),
    .ZN(_05677_));
 AOI22_X1 _22688_ (.A1(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .A2(_04550_),
    .B1(_04553_),
    .B2(\cs_registers_i.mhpmcounter[2][8] ),
    .ZN(_05678_));
 NOR2_X1 _22689_ (.A1(_04559_),
    .A2(_05678_),
    .ZN(_05679_));
 AOI22_X2 _22690_ (.A1(\cs_registers_i.dscratch0_q[8] ),
    .A2(_04511_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[8] ),
    .ZN(_05680_));
 AOI22_X2 _22691_ (.A1(net101),
    .A2(_04528_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .ZN(_05681_));
 INV_X1 _22692_ (.A(_01167_),
    .ZN(_05682_));
 AOI22_X2 _22693_ (.A1(_05682_),
    .A2(_05199_),
    .B1(net17),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .ZN(_05683_));
 NAND4_X2 _22694_ (.A1(_04247_),
    .A2(_05680_),
    .A3(_05681_),
    .A4(_05683_),
    .ZN(_05684_));
 NOR4_X4 _22695_ (.A1(_05675_),
    .A2(_05677_),
    .A3(_05679_),
    .A4(_05684_),
    .ZN(_05685_));
 AOI22_X4 _22696_ (.A1(_05672_),
    .A2(_05673_),
    .B1(_05685_),
    .B2(_04662_),
    .ZN(_05686_));
 AOI21_X4 _22697_ (.A(_05660_),
    .B1(_05686_),
    .B2(_04764_),
    .ZN(_05687_));
 CLKBUF_X3 _22698_ (.A(_05687_),
    .Z(_05688_));
 OAI21_X1 _22699_ (.A(_05654_),
    .B1(_05688_),
    .B2(_05465_),
    .ZN(_01205_));
 MUX2_X1 _22700_ (.A(_04912_),
    .B(_04913_),
    .S(_05513_),
    .Z(_05689_));
 MUX2_X1 _22701_ (.A(net68),
    .B(\load_store_unit_i.rdata_q[17] ),
    .S(_04911_),
    .Z(_05690_));
 MUX2_X1 _22702_ (.A(\load_store_unit_i.rdata_q[25] ),
    .B(net49),
    .S(_04911_),
    .Z(_05691_));
 MUX2_X1 _22703_ (.A(_05690_),
    .B(_05691_),
    .S(_05513_),
    .Z(_05692_));
 AOI22_X1 _22704_ (.A1(_04574_),
    .A2(_05689_),
    .B1(_05692_),
    .B2(_04581_),
    .ZN(_05693_));
 NAND2_X1 _22705_ (.A1(_04572_),
    .A2(_05693_),
    .ZN(_05694_));
 NAND2_X1 _22706_ (.A1(_04276_),
    .A2(_04459_),
    .ZN(_05695_));
 OR2_X1 _22707_ (.A1(_04455_),
    .A2(_05695_),
    .ZN(_05696_));
 OAI221_X1 _22708_ (.A(_04457_),
    .B1(_04308_),
    .B2(_04346_),
    .C1(_04307_),
    .C2(_04299_),
    .ZN(_05697_));
 NOR2_X1 _22709_ (.A1(_00563_),
    .A2(_04463_),
    .ZN(_05698_));
 NOR2_X1 _22710_ (.A1(_04625_),
    .A2(_04943_),
    .ZN(_05699_));
 NOR3_X2 _22711_ (.A1(_10493_),
    .A2(_05698_),
    .A3(_05699_),
    .ZN(_05700_));
 OAI21_X1 _22712_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B2(_11432_),
    .ZN(_05701_));
 AOI221_X1 _22713_ (.A(_04351_),
    .B1(_04358_),
    .B2(_15911_),
    .C1(_04362_),
    .C2(_15910_),
    .ZN(_05702_));
 AOI21_X1 _22714_ (.A(_05702_),
    .B1(_04353_),
    .B2(_15914_),
    .ZN(_05703_));
 AOI21_X1 _22715_ (.A(_05703_),
    .B1(_04369_),
    .B2(\alu_adder_result_ex[9] ),
    .ZN(_05704_));
 OAI221_X1 _22716_ (.A(_04393_),
    .B1(_05700_),
    .B2(_05701_),
    .C1(_05704_),
    .C2(_04390_),
    .ZN(_05705_));
 INV_X1 _22717_ (.A(_05705_),
    .ZN(_05706_));
 AND2_X1 _22718_ (.A1(_05697_),
    .A2(_05706_),
    .ZN(_05707_));
 BUF_X2 _22719_ (.A(\cs_registers_i.mhpmcounter[2][41] ),
    .Z(_05708_));
 AOI22_X2 _22720_ (.A1(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(_05708_),
    .ZN(_05709_));
 NOR2_X2 _22721_ (.A1(_04558_),
    .A2(_05709_),
    .ZN(_05710_));
 AOI22_X1 _22722_ (.A1(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\cs_registers_i.mhpmcounter[2][9] ),
    .ZN(_05711_));
 OR2_X1 _22723_ (.A1(_04559_),
    .A2(_05711_),
    .ZN(_05712_));
 AOI22_X2 _22724_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(_04521_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .ZN(_05713_));
 AOI222_X2 _22725_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(_04511_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .C1(_04775_),
    .C2(\cs_registers_i.dscratch1_q[9] ),
    .ZN(_05714_));
 OAI21_X2 _22726_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01168_),
    .ZN(_05715_));
 AOI221_X2 _22727_ (.A(_05715_),
    .B1(_04527_),
    .B2(net102),
    .C1(\cs_registers_i.mscratch_q[9] ),
    .C2(_04972_),
    .ZN(_05716_));
 NAND4_X2 _22728_ (.A1(_05712_),
    .A2(_05713_),
    .A3(_05714_),
    .A4(_05716_),
    .ZN(_05717_));
 NOR2_X4 _22729_ (.A1(_05710_),
    .A2(_05717_),
    .ZN(_05718_));
 AOI22_X4 _22730_ (.A1(_05696_),
    .A2(_05707_),
    .B1(_05718_),
    .B2(_04662_),
    .ZN(_05719_));
 MUX2_X2 _22731_ (.A(_05694_),
    .B(_05719_),
    .S(_04263_),
    .Z(_05720_));
 BUF_X2 _22732_ (.A(_05720_),
    .Z(_05721_));
 MUX2_X1 _22733_ (.A(_05721_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S(_05376_),
    .Z(_01206_));
 MUX2_X1 _22734_ (.A(_00564_),
    .B(_04997_),
    .S(_04463_),
    .Z(_05722_));
 NAND2_X1 _22735_ (.A1(_11432_),
    .A2(_05722_),
    .ZN(_05723_));
 INV_X1 _22736_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .ZN(_05724_));
 AOI21_X1 _22737_ (.A(_11406_),
    .B1(_05724_),
    .B2(_10310_),
    .ZN(_05725_));
 AOI21_X2 _22738_ (.A(_03493_),
    .B1(_05723_),
    .B2(_05725_),
    .ZN(_05726_));
 AOI22_X1 _22739_ (.A1(_15919_),
    .A2(_04358_),
    .B1(_04361_),
    .B2(_15918_),
    .ZN(_05727_));
 MUX2_X1 _22740_ (.A(_15922_),
    .B(_05727_),
    .S(_04664_),
    .Z(_05728_));
 AOI22_X1 _22741_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_04367_),
    .B1(_05475_),
    .B2(_04456_),
    .ZN(_05729_));
 NAND3_X1 _22742_ (.A1(_05726_),
    .A2(_05728_),
    .A3(_05729_),
    .ZN(_05730_));
 OAI21_X1 _22743_ (.A(_04281_),
    .B1(_04292_),
    .B2(_04990_),
    .ZN(_05731_));
 MUX2_X1 _22744_ (.A(_05122_),
    .B(_05130_),
    .S(_04452_),
    .Z(_05732_));
 OAI21_X1 _22745_ (.A(_05731_),
    .B1(_05732_),
    .B2(_04281_),
    .ZN(_05733_));
 AND2_X1 _22746_ (.A1(_04275_),
    .A2(_04459_),
    .ZN(_05734_));
 AOI221_X2 _22747_ (.A(_05730_),
    .B1(_05733_),
    .B2(_05734_),
    .C1(_05480_),
    .C2(_05009_),
    .ZN(_05735_));
 AOI22_X2 _22748_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(_04520_),
    .B1(_04542_),
    .B2(\cs_registers_i.csr_mepc_o[10] ),
    .ZN(_05736_));
 NAND2_X1 _22749_ (.A1(\cs_registers_i.mscratch_q[10] ),
    .A2(_04523_),
    .ZN(_05737_));
 AOI222_X2 _22750_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(net16),
    .B1(_04772_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C1(_04529_),
    .C2(\cs_registers_i.dscratch1_q[10] ),
    .ZN(_05738_));
 INV_X1 _22751_ (.A(_01169_),
    .ZN(_05739_));
 AOI221_X2 _22752_ (.A(_05231_),
    .B1(_05199_),
    .B2(_05739_),
    .C1(net72),
    .C2(_04526_),
    .ZN(_05740_));
 NAND4_X2 _22753_ (.A1(_05736_),
    .A2(_05737_),
    .A3(_05738_),
    .A4(_05740_),
    .ZN(_05741_));
 BUF_X2 _22754_ (.A(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .Z(_05742_));
 AOI22_X2 _22755_ (.A1(_05742_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(\cs_registers_i.mhpmcounter[2][42] ),
    .ZN(_05743_));
 INV_X1 _22756_ (.A(_05743_),
    .ZN(_05744_));
 NOR2_X4 _22757_ (.A1(_03551_),
    .A2(_04236_),
    .ZN(_05745_));
 OAI21_X1 _22758_ (.A(_03512_),
    .B1(_04234_),
    .B2(_15869_),
    .ZN(_05746_));
 NAND3_X1 _22759_ (.A1(_10922_),
    .A2(_03533_),
    .A3(_03514_),
    .ZN(_05747_));
 NOR2_X2 _22760_ (.A1(_05746_),
    .A2(_05747_),
    .ZN(_05748_));
 CLKBUF_X2 _22761_ (.A(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .Z(_05749_));
 BUF_X1 _22762_ (.A(\cs_registers_i.mhpmcounter[2][10] ),
    .Z(_05750_));
 AOI22_X1 _22763_ (.A1(_05749_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(_05750_),
    .ZN(_05751_));
 INV_X1 _22764_ (.A(_05751_),
    .ZN(_05752_));
 AOI221_X2 _22765_ (.A(_05741_),
    .B1(_05744_),
    .B2(_05745_),
    .C1(_05748_),
    .C2(_05752_),
    .ZN(_05753_));
 AOI221_X2 _22766_ (.A(_05735_),
    .B1(_05753_),
    .B2(_04662_),
    .C1(_04391_),
    .C2(_05726_),
    .ZN(_05754_));
 MUX2_X1 _22767_ (.A(_04979_),
    .B(_04980_),
    .S(_05513_),
    .Z(_05755_));
 MUX2_X1 _22768_ (.A(net39),
    .B(\load_store_unit_i.rdata_q[18] ),
    .S(_04911_),
    .Z(_05756_));
 MUX2_X1 _22769_ (.A(\load_store_unit_i.rdata_q[26] ),
    .B(net59),
    .S(_04911_),
    .Z(_05757_));
 MUX2_X1 _22770_ (.A(_05756_),
    .B(_05757_),
    .S(_05513_),
    .Z(_05758_));
 AOI22_X1 _22771_ (.A1(_04574_),
    .A2(_05755_),
    .B1(_05758_),
    .B2(_04582_),
    .ZN(_05759_));
 NAND2_X1 _22772_ (.A1(_04572_),
    .A2(_05759_),
    .ZN(_05760_));
 MUX2_X2 _22773_ (.A(_05754_),
    .B(_05760_),
    .S(_04906_),
    .Z(_05761_));
 CLKBUF_X2 _22774_ (.A(_05761_),
    .Z(_05762_));
 MUX2_X1 _22775_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .S(_05376_),
    .Z(_01207_));
 MUX2_X1 _22776_ (.A(net40),
    .B(\load_store_unit_i.rdata_q[19] ),
    .S(_04584_),
    .Z(_05763_));
 MUX2_X1 _22777_ (.A(\load_store_unit_i.rdata_q[27] ),
    .B(net62),
    .S(_04911_),
    .Z(_05764_));
 MUX2_X1 _22778_ (.A(_05763_),
    .B(_05764_),
    .S(_05513_),
    .Z(_05765_));
 MUX2_X1 _22779_ (.A(_04767_),
    .B(_04768_),
    .S(_04570_),
    .Z(_05766_));
 AOI22_X1 _22780_ (.A1(_04582_),
    .A2(_05765_),
    .B1(_05766_),
    .B2(_04574_),
    .ZN(_05767_));
 AND3_X1 _22781_ (.A1(_04611_),
    .A2(_04572_),
    .A3(_05767_),
    .ZN(_05768_));
 NOR2_X1 _22782_ (.A1(_00565_),
    .A2(_04502_),
    .ZN(_05769_));
 NOR2_X1 _22783_ (.A1(_05079_),
    .A2(_04810_),
    .ZN(_05770_));
 NOR3_X2 _22784_ (.A1(_10493_),
    .A2(_05769_),
    .A3(_05770_),
    .ZN(_05771_));
 OAI21_X1 _22785_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B2(_12102_),
    .ZN(_05772_));
 NOR2_X1 _22786_ (.A1(_05771_),
    .A2(_05772_),
    .ZN(_05773_));
 AOI221_X2 _22787_ (.A(_04351_),
    .B1(_04359_),
    .B2(_15927_),
    .C1(_04362_),
    .C2(_15926_),
    .ZN(_05774_));
 AOI21_X1 _22788_ (.A(_05774_),
    .B1(_04353_),
    .B2(_15930_),
    .ZN(_05775_));
 AOI21_X1 _22789_ (.A(_05775_),
    .B1(_04369_),
    .B2(\alu_adder_result_ex[11] ),
    .ZN(_05776_));
 AOI21_X1 _22790_ (.A(_04390_),
    .B1(_05476_),
    .B2(_05776_),
    .ZN(_05777_));
 NOR2_X1 _22791_ (.A1(_00550_),
    .A2(_04728_),
    .ZN(_05778_));
 AOI221_X2 _22792_ (.A(_05778_),
    .B1(_04738_),
    .B2(\cs_registers_i.mscratch_q[11] ),
    .C1(net135),
    .C2(_04742_),
    .ZN(_05779_));
 AOI221_X2 _22793_ (.A(_04741_),
    .B1(_04733_),
    .B2(\cs_registers_i.mie_q[15] ),
    .C1(net73),
    .C2(_04743_),
    .ZN(_05780_));
 AOI22_X2 _22794_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_04748_),
    .B1(_04749_),
    .B2(\cs_registers_i.dscratch1_q[11] ),
    .ZN(_05781_));
 AOI22_X2 _22795_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_04736_),
    .B1(_04747_),
    .B2(\cs_registers_i.mtval_q[11] ),
    .ZN(_05782_));
 NAND4_X2 _22796_ (.A1(_05779_),
    .A2(_05780_),
    .A3(_05781_),
    .A4(_05782_),
    .ZN(_05783_));
 AND4_X1 _22797_ (.A1(\cs_registers_i.mstack_d[0] ),
    .A2(_15507_),
    .A3(_03525_),
    .A4(_03553_),
    .ZN(_05784_));
 AOI221_X2 _22798_ (.A(_05784_),
    .B1(_05602_),
    .B2(\cs_registers_i.dcsr_q[11] ),
    .C1(\cs_registers_i.dscratch0_q[11] ),
    .C2(_04731_),
    .ZN(_05785_));
 CLKBUF_X2 _22799_ (.A(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .Z(_05786_));
 AOI22_X2 _22800_ (.A1(_05786_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(\cs_registers_i.mhpmcounter[2][43] ),
    .ZN(_05787_));
 OAI21_X1 _22801_ (.A(_05785_),
    .B1(_05787_),
    .B2(_04756_),
    .ZN(_05788_));
 BUF_X1 _22802_ (.A(\cs_registers_i.mhpmcounter[2][11] ),
    .Z(_05789_));
 AOI22_X1 _22803_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_04549_),
    .B1(_04552_),
    .B2(_05789_),
    .ZN(_05790_));
 NOR2_X1 _22804_ (.A1(_03532_),
    .A2(_05790_),
    .ZN(_05791_));
 OR3_X4 _22805_ (.A1(_05783_),
    .A2(_05788_),
    .A3(_05791_),
    .ZN(_05792_));
 AND3_X1 _22806_ (.A1(_04840_),
    .A2(_04722_),
    .A3(_04831_),
    .ZN(_05793_));
 OR4_X1 _22807_ (.A1(_05773_),
    .A2(_05777_),
    .A3(_05792_),
    .A4(_05793_),
    .ZN(_05794_));
 AOI21_X1 _22808_ (.A(_04458_),
    .B1(_04820_),
    .B2(_04720_),
    .ZN(_05795_));
 NOR2_X1 _22809_ (.A1(_04723_),
    .A2(_05795_),
    .ZN(_05796_));
 MUX2_X1 _22810_ (.A(_05054_),
    .B(_05049_),
    .S(_04453_),
    .Z(_05797_));
 AND2_X1 _22811_ (.A1(_04723_),
    .A2(_05797_),
    .ZN(_05798_));
 NOR3_X1 _22812_ (.A1(_04688_),
    .A2(_05796_),
    .A3(_05798_),
    .ZN(_05799_));
 NOR2_X2 _22813_ (.A1(_05794_),
    .A2(_05799_),
    .ZN(_05800_));
 AOI21_X4 _22814_ (.A(_05768_),
    .B1(_05800_),
    .B2(_04764_),
    .ZN(_05801_));
 BUF_X2 _22815_ (.A(_05801_),
    .Z(_05802_));
 MUX2_X1 _22816_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .S(_05376_),
    .Z(_01208_));
 CLKBUF_X3 _22817_ (.A(_04855_),
    .Z(_05803_));
 NAND2_X1 _22818_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .A2(_05803_),
    .ZN(_05804_));
 BUF_X4 _22819_ (.A(_05413_),
    .Z(_05805_));
 NAND2_X2 _22820_ (.A1(_04852_),
    .A2(_05805_),
    .ZN(_05806_));
 OAI21_X2 _22821_ (.A(_05804_),
    .B1(net445),
    .B2(_05806_),
    .ZN(_01209_));
 NAND2_X1 _22822_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .A2(_05416_),
    .ZN(_05807_));
 MUX2_X1 _22823_ (.A(_05038_),
    .B(_05039_),
    .S(_04596_),
    .Z(_05808_));
 MUX2_X1 _22824_ (.A(net41),
    .B(\load_store_unit_i.rdata_q[20] ),
    .S(_04593_),
    .Z(_05809_));
 MUX2_X1 _22825_ (.A(\load_store_unit_i.rdata_q[28] ),
    .B(net63),
    .S(_04593_),
    .Z(_05810_));
 MUX2_X1 _22826_ (.A(_05809_),
    .B(_05810_),
    .S(_05268_),
    .Z(_05811_));
 AOI22_X2 _22827_ (.A1(_04574_),
    .A2(_05808_),
    .B1(_05811_),
    .B2(_04582_),
    .ZN(_05812_));
 AOI21_X2 _22828_ (.A(_04600_),
    .B1(_04572_),
    .B2(_05812_),
    .ZN(_05813_));
 NAND2_X1 _22829_ (.A1(_00566_),
    .A2(_04625_),
    .ZN(_05814_));
 OAI21_X1 _22830_ (.A(_05814_),
    .B1(_05082_),
    .B2(_05079_),
    .ZN(_05815_));
 NAND2_X1 _22831_ (.A1(_12102_),
    .A2(_05815_),
    .ZN(_05816_));
 INV_X1 _22832_ (.A(_05816_),
    .ZN(_05817_));
 OAI21_X2 _22833_ (.A(_03449_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B2(_12102_),
    .ZN(_05818_));
 NAND2_X1 _22834_ (.A1(_04457_),
    .A2(_04723_),
    .ZN(_05819_));
 OAI221_X2 _22835_ (.A(_05661_),
    .B1(_05817_),
    .B2(_05818_),
    .C1(_05819_),
    .C2(_05055_),
    .ZN(_05820_));
 MUX2_X1 _22836_ (.A(_15935_),
    .B(_15934_),
    .S(_04363_),
    .Z(_05821_));
 NAND2_X1 _22837_ (.A1(_04665_),
    .A2(_05821_),
    .ZN(_05822_));
 OAI21_X1 _22838_ (.A(_05822_),
    .B1(_04665_),
    .B2(_15938_),
    .ZN(_05823_));
 AOI22_X2 _22839_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_04825_),
    .B1(_05823_),
    .B2(_05562_),
    .ZN(_05824_));
 AOI22_X1 _22840_ (.A1(_04707_),
    .A2(_04699_),
    .B1(_04828_),
    .B2(_04692_),
    .ZN(_05825_));
 NAND2_X1 _22841_ (.A1(_04702_),
    .A2(_04704_),
    .ZN(_05826_));
 MUX2_X1 _22842_ (.A(_05826_),
    .B(_04711_),
    .S(_04707_),
    .Z(_05827_));
 MUX2_X1 _22843_ (.A(_05825_),
    .B(_05827_),
    .S(_04720_),
    .Z(_05828_));
 INV_X1 _22844_ (.A(_05120_),
    .ZN(_05829_));
 MUX2_X1 _22845_ (.A(_04674_),
    .B(_04830_),
    .S(_04720_),
    .Z(_05830_));
 NAND2_X1 _22846_ (.A1(_04308_),
    .A2(_04276_),
    .ZN(_05831_));
 OAI221_X1 _22847_ (.A(_05824_),
    .B1(_05828_),
    .B2(_05829_),
    .C1(_05830_),
    .C2(_05831_),
    .ZN(_05832_));
 AOI21_X1 _22848_ (.A(_05820_),
    .B1(_05832_),
    .B2(_04815_),
    .ZN(_05833_));
 AOI22_X1 _22849_ (.A1(\cs_registers_i.mscratch_q[12] ),
    .A2(_04972_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[12] ),
    .ZN(_05834_));
 NAND2_X1 _22850_ (.A1(\cs_registers_i.mtval_q[12] ),
    .A2(_04520_),
    .ZN(_05835_));
 AND3_X1 _22851_ (.A1(_04247_),
    .A2(_05834_),
    .A3(_05835_),
    .ZN(_05836_));
 AOI222_X2 _22852_ (.A1(\cs_registers_i.dscratch1_q[12] ),
    .A2(_04775_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .C1(_05487_),
    .C2(\cs_registers_i.mstack_d[1] ),
    .ZN(_05837_));
 AOI22_X1 _22853_ (.A1(net74),
    .A2(_05490_),
    .B1(net17),
    .B2(\cs_registers_i.dcsr_q[12] ),
    .ZN(_05838_));
 NAND3_X1 _22854_ (.A1(_03501_),
    .A2(_15873_),
    .A3(_03542_),
    .ZN(_05839_));
 NOR3_X2 _22855_ (.A1(_03563_),
    .A2(_04512_),
    .A3(_05839_),
    .ZN(_05840_));
 INV_X1 _22856_ (.A(_00549_),
    .ZN(_05841_));
 AOI22_X1 _22857_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_04771_),
    .B1(_05840_),
    .B2(_05841_),
    .ZN(_05842_));
 AND4_X1 _22858_ (.A1(_05836_),
    .A2(_05837_),
    .A3(_05838_),
    .A4(_05842_),
    .ZN(_05843_));
 AOI22_X2 _22859_ (.A1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][44] ),
    .ZN(_05844_));
 AOI22_X2 _22860_ (.A1(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][12] ),
    .ZN(_05845_));
 OAI221_X2 _22861_ (.A(_05843_),
    .B1(_05844_),
    .B2(_05031_),
    .C1(_04560_),
    .C2(_05845_),
    .ZN(_05846_));
 NOR2_X2 _22862_ (.A1(_04563_),
    .A2(_05846_),
    .ZN(_05847_));
 NOR3_X2 _22863_ (.A1(_04906_),
    .A2(_05833_),
    .A3(_05847_),
    .ZN(_05848_));
 NOR2_X2 _22864_ (.A1(_05813_),
    .A2(_05848_),
    .ZN(_05849_));
 CLKBUF_X3 _22865_ (.A(_05849_),
    .Z(_05850_));
 OAI21_X1 _22866_ (.A(_05807_),
    .B1(_05850_),
    .B2(_05465_),
    .ZN(_01210_));
 MUX2_X1 _22867_ (.A(_05096_),
    .B(_05097_),
    .S(_05513_),
    .Z(_05851_));
 MUX2_X1 _22868_ (.A(net42),
    .B(\load_store_unit_i.rdata_q[21] ),
    .S(_04585_),
    .Z(_05852_));
 MUX2_X1 _22869_ (.A(\load_store_unit_i.rdata_q[29] ),
    .B(net64),
    .S(_04585_),
    .Z(_05853_));
 MUX2_X1 _22870_ (.A(_05852_),
    .B(_05853_),
    .S(_05513_),
    .Z(_05854_));
 AOI22_X2 _22871_ (.A1(_04574_),
    .A2(_05851_),
    .B1(_05854_),
    .B2(_04582_),
    .ZN(_05855_));
 NAND2_X1 _22872_ (.A1(_04572_),
    .A2(_05855_),
    .ZN(_05856_));
 NAND2_X1 _22873_ (.A1(_04611_),
    .A2(_05856_),
    .ZN(_05857_));
 NOR2_X2 _22874_ (.A1(_10310_),
    .A2(_04623_),
    .ZN(_05858_));
 NAND2_X1 _22875_ (.A1(_05104_),
    .A2(_05858_),
    .ZN(_05859_));
 OAI21_X2 _22876_ (.A(_05859_),
    .B1(_05858_),
    .B2(_04023_),
    .ZN(_05860_));
 INV_X1 _22877_ (.A(_15946_),
    .ZN(_05861_));
 AOI22_X1 _22878_ (.A1(_05861_),
    .A2(_04351_),
    .B1(_04367_),
    .B2(\alu_adder_result_ex[13] ),
    .ZN(_05862_));
 AOI22_X1 _22879_ (.A1(_15943_),
    .A2(_04359_),
    .B1(_04362_),
    .B2(_15942_),
    .ZN(_05863_));
 OAI21_X1 _22880_ (.A(_05862_),
    .B1(_05863_),
    .B2(_04351_),
    .ZN(_05864_));
 AOI221_X2 _22881_ (.A(_03493_),
    .B1(_11401_),
    .B2(_05860_),
    .C1(_05864_),
    .C2(_04814_),
    .ZN(_05865_));
 INV_X1 _22882_ (.A(_05865_),
    .ZN(_05866_));
 MUX2_X1 _22883_ (.A(_05008_),
    .B(_05010_),
    .S(_04453_),
    .Z(_05867_));
 NOR2_X1 _22884_ (.A1(_04412_),
    .A2(_04687_),
    .ZN(_05868_));
 AOI221_X2 _22885_ (.A(_05866_),
    .B1(_05867_),
    .B2(_05120_),
    .C1(_05119_),
    .C2(_05868_),
    .ZN(_05869_));
 NAND3_X1 _22886_ (.A1(_04410_),
    .A2(_04916_),
    .A3(_04917_),
    .ZN(_05870_));
 OAI21_X1 _22887_ (.A(_05870_),
    .B1(_04331_),
    .B2(_04431_),
    .ZN(_05871_));
 MUX2_X1 _22888_ (.A(_04990_),
    .B(_05871_),
    .S(_04453_),
    .Z(_05872_));
 AOI21_X1 _22889_ (.A(_05475_),
    .B1(_05872_),
    .B2(_04723_),
    .ZN(_05873_));
 OAI21_X2 _22890_ (.A(_05869_),
    .B1(_05873_),
    .B2(_04725_),
    .ZN(_05874_));
 CLKBUF_X3 _22891_ (.A(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .Z(_05875_));
 AOI22_X2 _22892_ (.A1(_05875_),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][45] ),
    .ZN(_05876_));
 NOR2_X1 _22893_ (.A1(_04558_),
    .A2(_05876_),
    .ZN(_05877_));
 CLKBUF_X2 _22894_ (.A(\cs_registers_i.mhpmcounter[2][13] ),
    .Z(_05878_));
 AOI22_X1 _22895_ (.A1(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(_05878_),
    .ZN(_05879_));
 NOR2_X1 _22896_ (.A1(_04783_),
    .A2(_05879_),
    .ZN(_05880_));
 AOI22_X1 _22897_ (.A1(\cs_registers_i.mscratch_q[13] ),
    .A2(_04524_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[13] ),
    .ZN(_05881_));
 AOI22_X2 _22898_ (.A1(\cs_registers_i.dscratch1_q[13] ),
    .A2(_04530_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[13] ),
    .ZN(_05882_));
 AOI22_X2 _22899_ (.A1(net75),
    .A2(_04528_),
    .B1(net17),
    .B2(\cs_registers_i.dcsr_q[13] ),
    .ZN(_05883_));
 OAI21_X1 _22900_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01170_),
    .ZN(_05884_));
 AOI221_X2 _22901_ (.A(_05884_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .C1(\cs_registers_i.dscratch0_q[13] ),
    .C2(_04771_),
    .ZN(_05885_));
 NAND4_X2 _22902_ (.A1(_05881_),
    .A2(_05882_),
    .A3(_05883_),
    .A4(_05885_),
    .ZN(_05886_));
 OR3_X2 _22903_ (.A1(_05877_),
    .A2(_05880_),
    .A3(_05886_),
    .ZN(_05887_));
 OAI21_X2 _22904_ (.A(_05874_),
    .B1(_05887_),
    .B2(_04563_),
    .ZN(_05888_));
 OAI21_X4 _22905_ (.A(_05857_),
    .B1(_05888_),
    .B2(_04906_),
    .ZN(_05889_));
 BUF_X2 _22906_ (.A(_05889_),
    .Z(_05890_));
 MUX2_X1 _22907_ (.A(_05890_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .S(_05376_),
    .Z(_01211_));
 MUX2_X1 _22908_ (.A(net43),
    .B(\load_store_unit_i.rdata_q[22] ),
    .S(_04584_),
    .Z(_05891_));
 MUX2_X1 _22909_ (.A(\load_store_unit_i.rdata_q[30] ),
    .B(net65),
    .S(_04911_),
    .Z(_05892_));
 MUX2_X1 _22910_ (.A(_05891_),
    .B(_05892_),
    .S(_04570_),
    .Z(_05893_));
 MUX2_X1 _22911_ (.A(_05206_),
    .B(_05207_),
    .S(_04570_),
    .Z(_05894_));
 AOI22_X1 _22912_ (.A1(_04582_),
    .A2(_05893_),
    .B1(_05894_),
    .B2(_04574_),
    .ZN(_05895_));
 AND3_X1 _22913_ (.A1(_04905_),
    .A2(_04572_),
    .A3(_05895_),
    .ZN(_05896_));
 NOR2_X1 _22914_ (.A1(_04026_),
    .A2(_05858_),
    .ZN(_05897_));
 AOI21_X1 _22915_ (.A(_05897_),
    .B1(_05858_),
    .B2(_05158_),
    .ZN(_05898_));
 NOR2_X2 _22916_ (.A1(_11407_),
    .A2(_05898_),
    .ZN(_05899_));
 NOR3_X1 _22917_ (.A1(_04725_),
    .A2(_04411_),
    .A3(_04670_),
    .ZN(_05900_));
 AND3_X1 _22918_ (.A1(_04457_),
    .A2(_04685_),
    .A3(_04432_),
    .ZN(_05901_));
 NOR4_X2 _22919_ (.A1(_05477_),
    .A2(_05899_),
    .A3(_05900_),
    .A4(_05901_),
    .ZN(_05902_));
 OR3_X1 _22920_ (.A1(_04293_),
    .A2(_04298_),
    .A3(_04928_),
    .ZN(_05903_));
 OAI21_X1 _22921_ (.A(_04307_),
    .B1(_04298_),
    .B2(_04293_),
    .ZN(_05904_));
 AOI21_X1 _22922_ (.A(_04722_),
    .B1(_05903_),
    .B2(_05904_),
    .ZN(_05905_));
 AOI21_X1 _22923_ (.A(_04308_),
    .B1(_04720_),
    .B2(_04924_),
    .ZN(_05906_));
 OR2_X1 _22924_ (.A1(_04340_),
    .A2(_04720_),
    .ZN(_05907_));
 AOI21_X2 _22925_ (.A(_05905_),
    .B1(_05906_),
    .B2(_05907_),
    .ZN(_05908_));
 MUX2_X1 _22926_ (.A(_15951_),
    .B(_15950_),
    .S(_04363_),
    .Z(_05909_));
 NAND2_X1 _22927_ (.A1(_04665_),
    .A2(_05909_),
    .ZN(_05910_));
 OAI21_X1 _22928_ (.A(_05910_),
    .B1(_04665_),
    .B2(_15954_),
    .ZN(_05911_));
 AOI22_X2 _22929_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_04825_),
    .B1(_05911_),
    .B2(_05562_),
    .ZN(_05912_));
 OAI221_X2 _22930_ (.A(_05902_),
    .B1(_05908_),
    .B2(_04688_),
    .C1(_05912_),
    .C2(_04391_),
    .ZN(_05913_));
 CLKBUF_X3 _22931_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .Z(_05914_));
 AOI22_X4 _22932_ (.A1(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(_05914_),
    .ZN(_05915_));
 NOR2_X2 _22933_ (.A1(_05031_),
    .A2(_05915_),
    .ZN(_05916_));
 AOI22_X1 _22934_ (.A1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][14] ),
    .ZN(_05917_));
 NOR2_X1 _22935_ (.A1(_04783_),
    .A2(_05917_),
    .ZN(_05918_));
 AOI22_X1 _22936_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(_04521_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .ZN(_05919_));
 AOI222_X2 _22937_ (.A1(\cs_registers_i.dscratch0_q[14] ),
    .A2(_04511_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[14] ),
    .C1(_04775_),
    .C2(\cs_registers_i.dscratch1_q[14] ),
    .ZN(_05920_));
 OAI21_X1 _22938_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01171_),
    .ZN(_05921_));
 AOI221_X2 _22939_ (.A(_05921_),
    .B1(_04527_),
    .B2(net76),
    .C1(\cs_registers_i.mscratch_q[14] ),
    .C2(_04972_),
    .ZN(_05922_));
 NAND3_X2 _22940_ (.A1(_05919_),
    .A2(_05920_),
    .A3(_05922_),
    .ZN(_05923_));
 NOR3_X4 _22941_ (.A1(_05916_),
    .A2(_05918_),
    .A3(_05923_),
    .ZN(_05924_));
 INV_X1 _22942_ (.A(_05924_),
    .ZN(_05925_));
 OAI21_X2 _22943_ (.A(_05913_),
    .B1(_05925_),
    .B2(_04563_),
    .ZN(_05926_));
 AOI21_X4 _22944_ (.A(_05896_),
    .B1(_05926_),
    .B2(_04600_),
    .ZN(_05927_));
 BUF_X2 _22945_ (.A(_05927_),
    .Z(_05928_));
 BUF_X4 _22946_ (.A(_05375_),
    .Z(_05929_));
 MUX2_X1 _22947_ (.A(_05928_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .S(_05929_),
    .Z(_01212_));
 NAND3_X1 _22948_ (.A1(_05513_),
    .A2(_04589_),
    .A3(net61),
    .ZN(_05930_));
 NAND3_X1 _22949_ (.A1(_04577_),
    .A2(_04586_),
    .A3(_04568_),
    .ZN(_05931_));
 AOI21_X1 _22950_ (.A(_05271_),
    .B1(_05930_),
    .B2(_05931_),
    .ZN(_05932_));
 AND3_X1 _22951_ (.A1(_04577_),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .A3(_04581_),
    .ZN(_05933_));
 OAI21_X1 _22952_ (.A(_04594_),
    .B1(_05932_),
    .B2(_05933_),
    .ZN(_05934_));
 AND3_X1 _22953_ (.A1(_05268_),
    .A2(_04586_),
    .A3(net66),
    .ZN(_05935_));
 AND3_X1 _22954_ (.A1(_04577_),
    .A2(_04589_),
    .A3(net44),
    .ZN(_05936_));
 OAI21_X1 _22955_ (.A(_05272_),
    .B1(_05935_),
    .B2(_05936_),
    .ZN(_05937_));
 AND3_X1 _22956_ (.A1(_04589_),
    .A2(\load_store_unit_i.rdata_q[31] ),
    .A3(_04581_),
    .ZN(_05938_));
 OAI21_X1 _22957_ (.A(_05421_),
    .B1(_05932_),
    .B2(_05938_),
    .ZN(_05939_));
 NAND4_X2 _22958_ (.A1(_04572_),
    .A2(_05934_),
    .A3(_05937_),
    .A4(_05939_),
    .ZN(_05940_));
 INV_X1 _22959_ (.A(_15958_),
    .ZN(_05941_));
 AOI22_X1 _22960_ (.A1(_05941_),
    .A2(_04352_),
    .B1(_04367_),
    .B2(\alu_adder_result_ex[15] ),
    .ZN(_05942_));
 AOI22_X1 _22961_ (.A1(_15959_),
    .A2(_04360_),
    .B1(_04983_),
    .B2(_15962_),
    .ZN(_05943_));
 OAI21_X1 _22962_ (.A(_05942_),
    .B1(_05943_),
    .B2(_04353_),
    .ZN(_05944_));
 NAND2_X1 _22963_ (.A1(_04814_),
    .A2(_05944_),
    .ZN(_05945_));
 MUX2_X1 _22964_ (.A(_00659_),
    .B(_05219_),
    .S(_05858_),
    .Z(_05946_));
 OR2_X2 _22965_ (.A1(_11407_),
    .A2(_05946_),
    .ZN(_05947_));
 AND3_X2 _22966_ (.A1(_05661_),
    .A2(_05945_),
    .A3(_05947_),
    .ZN(_05948_));
 NAND2_X1 _22967_ (.A1(_04840_),
    .A2(_04722_),
    .ZN(_05949_));
 NAND2_X1 _22968_ (.A1(_04429_),
    .A2(_04326_),
    .ZN(_05950_));
 NOR2_X1 _22969_ (.A1(_04431_),
    .A2(_04698_),
    .ZN(_05951_));
 AOI22_X1 _22970_ (.A1(_05950_),
    .A2(_05951_),
    .B1(_04705_),
    .B2(_04707_),
    .ZN(_05952_));
 MUX2_X1 _22971_ (.A(_04695_),
    .B(_05952_),
    .S(_04453_),
    .Z(_05953_));
 NOR2_X1 _22972_ (.A1(_04399_),
    .A2(_04675_),
    .ZN(_05954_));
 NOR2_X1 _22973_ (.A1(_04333_),
    .A2(_04292_),
    .ZN(_05955_));
 AOI21_X1 _22974_ (.A(_04307_),
    .B1(_05954_),
    .B2(_05955_),
    .ZN(_05956_));
 OAI221_X1 _22975_ (.A(_05948_),
    .B1(_05949_),
    .B2(_05953_),
    .C1(_05831_),
    .C2(_05956_),
    .ZN(_05957_));
 MUX2_X1 _22976_ (.A(_04684_),
    .B(_04883_),
    .S(_04720_),
    .Z(_05958_));
 AOI21_X2 _22977_ (.A(_05957_),
    .B1(_05958_),
    .B2(_05120_),
    .ZN(_05959_));
 AOI22_X1 _22978_ (.A1(\cs_registers_i.mscratch_q[15] ),
    .A2(_04524_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[15] ),
    .ZN(_05960_));
 AOI22_X1 _22979_ (.A1(\cs_registers_i.dscratch1_q[15] ),
    .A2(_04775_),
    .B1(net17),
    .B2(\cs_registers_i.dcsr_q[15] ),
    .ZN(_05961_));
 AOI22_X1 _22980_ (.A1(net77),
    .A2(_04528_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[15] ),
    .ZN(_05962_));
 OAI21_X1 _22981_ (.A(_04533_),
    .B1(_04536_),
    .B2(_01172_),
    .ZN(_05963_));
 AOI221_X2 _22982_ (.A(_05963_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .C1(\cs_registers_i.dscratch0_q[15] ),
    .C2(net16),
    .ZN(_05964_));
 AND4_X1 _22983_ (.A1(_05960_),
    .A2(_05961_),
    .A3(_05962_),
    .A4(_05964_),
    .ZN(_05965_));
 BUF_X2 _22984_ (.A(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .Z(_05966_));
 BUF_X2 _22985_ (.A(\cs_registers_i.mhpmcounter[2][47] ),
    .Z(_05967_));
 AOI22_X4 _22986_ (.A1(_05966_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(_05967_),
    .ZN(_05968_));
 AOI22_X2 _22987_ (.A1(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][15] ),
    .ZN(_05969_));
 OAI221_X2 _22988_ (.A(_05965_),
    .B1(_05968_),
    .B2(_04557_),
    .C1(_04783_),
    .C2(_05969_),
    .ZN(_05970_));
 NOR2_X1 _22989_ (.A1(_04393_),
    .A2(_05970_),
    .ZN(_05971_));
 NOR2_X1 _22990_ (.A1(_05959_),
    .A2(_05971_),
    .ZN(_05972_));
 MUX2_X2 _22991_ (.A(_05940_),
    .B(_05972_),
    .S(_04263_),
    .Z(_05973_));
 BUF_X4 _22992_ (.A(_05973_),
    .Z(_05974_));
 MUX2_X1 _22993_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .S(_05929_),
    .Z(_01213_));
 NAND2_X1 _22994_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .A2(_05416_),
    .ZN(_05975_));
 MUX2_X1 _22995_ (.A(net38),
    .B(net67),
    .S(_04593_),
    .Z(_05976_));
 NAND2_X1 _22996_ (.A1(_04596_),
    .A2(_05976_),
    .ZN(_05977_));
 AOI21_X1 _22997_ (.A(_05263_),
    .B1(\load_store_unit_i.rdata_q[24] ),
    .B2(_04594_),
    .ZN(_05978_));
 OAI21_X1 _22998_ (.A(_05977_),
    .B1(_05978_),
    .B2(_05421_),
    .ZN(_05979_));
 AOI21_X1 _22999_ (.A(_04580_),
    .B1(_04582_),
    .B2(_05979_),
    .ZN(_05980_));
 NOR2_X2 _23000_ (.A1(_04600_),
    .A2(_05980_),
    .ZN(_05981_));
 NAND2_X1 _23001_ (.A1(_04308_),
    .A2(_04307_),
    .ZN(_05982_));
 OAI21_X1 _23002_ (.A(_05982_),
    .B1(_05953_),
    .B2(_04308_),
    .ZN(_05983_));
 NAND2_X1 _23003_ (.A1(_04276_),
    .A2(_05983_),
    .ZN(_05984_));
 NAND2_X1 _23004_ (.A1(_15553_),
    .A2(_04624_),
    .ZN(_05985_));
 NOR2_X1 _23005_ (.A1(_04490_),
    .A2(_04474_),
    .ZN(_05986_));
 AOI21_X1 _23006_ (.A(_05986_),
    .B1(_04492_),
    .B2(_04639_),
    .ZN(_05987_));
 AOI21_X2 _23007_ (.A(_15725_),
    .B1(_05987_),
    .B2(_15726_),
    .ZN(_05988_));
 XNOR2_X2 _23008_ (.A(_15730_),
    .B(_05988_),
    .ZN(_05989_));
 NAND2_X1 _23009_ (.A1(_04463_),
    .A2(_05989_),
    .ZN(_05990_));
 NAND3_X2 _23010_ (.A1(_11432_),
    .A2(_05985_),
    .A3(_05990_),
    .ZN(_05991_));
 AOI21_X1 _23011_ (.A(_11406_),
    .B1(_03670_),
    .B2(_10310_),
    .ZN(_05992_));
 AOI21_X2 _23012_ (.A(_04662_),
    .B1(_05991_),
    .B2(_05992_),
    .ZN(_05993_));
 AOI221_X1 _23013_ (.A(_04351_),
    .B1(_04358_),
    .B2(_15967_),
    .C1(_04362_),
    .C2(_15966_),
    .ZN(_05994_));
 AOI21_X1 _23014_ (.A(_05994_),
    .B1(_04353_),
    .B2(_15970_),
    .ZN(_05995_));
 AOI21_X1 _23015_ (.A(_05995_),
    .B1(_04368_),
    .B2(\alu_adder_result_ex[16] ),
    .ZN(_05996_));
 OAI21_X2 _23016_ (.A(_05993_),
    .B1(_05996_),
    .B2(_04390_),
    .ZN(_05997_));
 NOR2_X1 _23017_ (.A1(_04725_),
    .A2(_04722_),
    .ZN(_05998_));
 MUX2_X1 _23018_ (.A(_04307_),
    .B(_04676_),
    .S(_05955_),
    .Z(_05999_));
 NOR2_X1 _23019_ (.A1(_04725_),
    .A2(_04308_),
    .ZN(_06000_));
 AOI221_X2 _23020_ (.A(_05997_),
    .B1(_05998_),
    .B2(_05999_),
    .C1(_05958_),
    .C2(_06000_),
    .ZN(_06001_));
 AOI22_X2 _23021_ (.A1(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][48] ),
    .ZN(_06002_));
 NOR2_X1 _23022_ (.A1(_04558_),
    .A2(_06002_),
    .ZN(_06003_));
 BUF_X2 _23023_ (.A(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .Z(_06004_));
 AOI22_X2 _23024_ (.A1(_06004_),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][16] ),
    .ZN(_06005_));
 NOR2_X2 _23025_ (.A1(_04560_),
    .A2(_06005_),
    .ZN(_06006_));
 AOI22_X2 _23026_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(_04515_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .ZN(_06007_));
 AOI22_X4 _23027_ (.A1(\cs_registers_i.dscratch0_q[16] ),
    .A2(_04511_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[16] ),
    .ZN(_06008_));
 AOI222_X2 _23028_ (.A1(net136),
    .A2(_04518_),
    .B1(_05022_),
    .B2(\cs_registers_i.mtval_q[16] ),
    .C1(\cs_registers_i.mscratch_q[16] ),
    .C2(_04524_),
    .ZN(_06009_));
 OAI21_X1 _23029_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01173_),
    .ZN(_06010_));
 AOI221_X2 _23030_ (.A(_06010_),
    .B1(_04527_),
    .B2(net78),
    .C1(\cs_registers_i.csr_mepc_o[16] ),
    .C2(_05074_),
    .ZN(_06011_));
 NAND4_X4 _23031_ (.A1(_06007_),
    .A2(_06008_),
    .A3(_06009_),
    .A4(_06011_),
    .ZN(_06012_));
 NOR3_X4 _23032_ (.A1(_06003_),
    .A2(_06006_),
    .A3(_06012_),
    .ZN(_06013_));
 AOI22_X4 _23033_ (.A1(_05984_),
    .A2(_06001_),
    .B1(_06013_),
    .B2(_04662_),
    .ZN(_06014_));
 AOI21_X4 _23034_ (.A(_05981_),
    .B1(_06014_),
    .B2(_04764_),
    .ZN(_06015_));
 CLKBUF_X3 _23035_ (.A(_06015_),
    .Z(_06016_));
 OAI21_X1 _23036_ (.A(_05975_),
    .B1(_06016_),
    .B2(_05465_),
    .ZN(_01214_));
 NAND3_X1 _23037_ (.A1(_05421_),
    .A2(_05378_),
    .A3(_05383_),
    .ZN(_06017_));
 MUX2_X1 _23038_ (.A(net46),
    .B(\load_store_unit_i.rdata_q[25] ),
    .S(_04586_),
    .Z(_06018_));
 OAI21_X1 _23039_ (.A(_06017_),
    .B1(_06018_),
    .B2(_05421_),
    .ZN(_06019_));
 INV_X1 _23040_ (.A(_06019_),
    .ZN(_06020_));
 AOI21_X4 _23041_ (.A(_04617_),
    .B1(_06020_),
    .B2(_04583_),
    .ZN(_06021_));
 AOI21_X1 _23042_ (.A(_10310_),
    .B1(_15556_),
    .B2(_04625_),
    .ZN(_06022_));
 NAND2_X1 _23043_ (.A1(_04640_),
    .A2(_04642_),
    .ZN(_06023_));
 NAND3_X1 _23044_ (.A1(_15700_),
    .A2(_04640_),
    .A3(_04652_),
    .ZN(_06024_));
 NAND3_X2 _23045_ (.A1(_04495_),
    .A2(_06023_),
    .A3(_06024_),
    .ZN(_06025_));
 XNOR2_X2 _23046_ (.A(_04472_),
    .B(_06025_),
    .ZN(_06026_));
 OAI21_X2 _23047_ (.A(_06022_),
    .B1(_06026_),
    .B2(_04626_),
    .ZN(_06027_));
 AOI21_X1 _23048_ (.A(_11407_),
    .B1(_03800_),
    .B2(net300),
    .ZN(_06028_));
 NAND2_X1 _23049_ (.A1(_06027_),
    .A2(_06028_),
    .ZN(_06029_));
 AOI221_X1 _23050_ (.A(_04351_),
    .B1(_04359_),
    .B2(_15975_),
    .C1(_04983_),
    .C2(_15974_),
    .ZN(_06030_));
 AOI21_X1 _23051_ (.A(_06030_),
    .B1(_04370_),
    .B2(_15978_),
    .ZN(_06031_));
 AOI21_X1 _23052_ (.A(_06031_),
    .B1(_04825_),
    .B2(\alu_adder_result_ex[17] ),
    .ZN(_06032_));
 OAI21_X1 _23053_ (.A(_06029_),
    .B1(_06032_),
    .B2(_04390_),
    .ZN(_06033_));
 CLKBUF_X3 _23054_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .Z(_06034_));
 AOI22_X2 _23055_ (.A1(_06034_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(\cs_registers_i.mhpmcounter[2][49] ),
    .ZN(_06035_));
 NOR3_X1 _23056_ (.A1(_03551_),
    .A2(_04236_),
    .A3(_06035_),
    .ZN(_06036_));
 BUF_X2 _23057_ (.A(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .Z(_06037_));
 BUF_X2 _23058_ (.A(\cs_registers_i.mhpmcounter[2][17] ),
    .Z(_06038_));
 AOI22_X2 _23059_ (.A1(_06037_),
    .A2(_04549_),
    .B1(_04552_),
    .B2(_06038_),
    .ZN(_06039_));
 NOR2_X1 _23060_ (.A1(_04559_),
    .A2(_06039_),
    .ZN(_06040_));
 AOI22_X1 _23061_ (.A1(net142),
    .A2(_04517_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[17] ),
    .ZN(_06041_));
 AOI22_X1 _23062_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(_04972_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[17] ),
    .ZN(_06042_));
 NAND2_X1 _23063_ (.A1(_06041_),
    .A2(_06042_),
    .ZN(_06043_));
 AND2_X1 _23064_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(_04514_),
    .ZN(_06044_));
 INV_X1 _23065_ (.A(\cs_registers_i.dscratch0_q[17] ),
    .ZN(_06045_));
 INV_X1 _23066_ (.A(\cs_registers_i.mstatus_q[1] ),
    .ZN(_06046_));
 OAI33_X1 _23067_ (.A1(_06045_),
    .A2(_04509_),
    .A3(_04730_),
    .B1(_05452_),
    .B2(_11072_),
    .B3(_06046_),
    .ZN(_06047_));
 INV_X1 _23068_ (.A(\cs_registers_i.dscratch1_q[17] ),
    .ZN(_06048_));
 OAI221_X1 _23069_ (.A(_04533_),
    .B1(_04536_),
    .B2(_01174_),
    .C1(_05450_),
    .C2(_06048_),
    .ZN(_06049_));
 INV_X1 _23070_ (.A(net79),
    .ZN(_06050_));
 INV_X1 _23071_ (.A(\cs_registers_i.csr_depc_o[17] ),
    .ZN(_06051_));
 OAI22_X1 _23072_ (.A1(_06050_),
    .A2(_04256_),
    .B1(_04539_),
    .B2(_06051_),
    .ZN(_06052_));
 OR4_X2 _23073_ (.A1(_06044_),
    .A2(_06047_),
    .A3(_06049_),
    .A4(_06052_),
    .ZN(_06053_));
 OR4_X4 _23074_ (.A1(_06036_),
    .A2(_06040_),
    .A3(_06043_),
    .A4(_06053_),
    .ZN(_06054_));
 NOR2_X1 _23075_ (.A1(_06033_),
    .A2(_06054_),
    .ZN(_06055_));
 OAI21_X2 _23076_ (.A(_06055_),
    .B1(_05908_),
    .B2(_04342_),
    .ZN(_06056_));
 AOI21_X1 _23077_ (.A(_05177_),
    .B1(_04411_),
    .B2(_04293_),
    .ZN(_06057_));
 NAND2_X1 _23078_ (.A1(_04723_),
    .A2(_06057_),
    .ZN(_06058_));
 AOI21_X2 _23079_ (.A(_04688_),
    .B1(_05982_),
    .B2(_06058_),
    .ZN(_06059_));
 NOR3_X4 _23080_ (.A1(_04906_),
    .A2(_06056_),
    .A3(_06059_),
    .ZN(_06060_));
 NOR2_X4 _23081_ (.A1(_06021_),
    .A2(_06060_),
    .ZN(_06061_));
 BUF_X2 _23082_ (.A(_06061_),
    .Z(_06062_));
 MUX2_X1 _23083_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .S(_05929_),
    .Z(_01215_));
 NAND3_X1 _23084_ (.A1(_04596_),
    .A2(_05423_),
    .A3(_05419_),
    .ZN(_06063_));
 MUX2_X1 _23085_ (.A(net47),
    .B(\load_store_unit_i.rdata_q[26] ),
    .S(_04586_),
    .Z(_06064_));
 OAI21_X1 _23086_ (.A(_06063_),
    .B1(_06064_),
    .B2(_05421_),
    .ZN(_06065_));
 INV_X1 _23087_ (.A(_06065_),
    .ZN(_06066_));
 AOI21_X4 _23088_ (.A(_04617_),
    .B1(_06066_),
    .B2(_04583_),
    .ZN(_06067_));
 AOI22_X1 _23089_ (.A1(_15983_),
    .A2(_04359_),
    .B1(_04983_),
    .B2(_15986_),
    .ZN(_06068_));
 MUX2_X1 _23090_ (.A(_15982_),
    .B(_06068_),
    .S(_04664_),
    .Z(_06069_));
 NAND2_X1 _23091_ (.A1(_05116_),
    .A2(_06069_),
    .ZN(_06070_));
 AOI221_X1 _23092_ (.A(_06070_),
    .B1(_05872_),
    .B2(_05120_),
    .C1(net450),
    .C2(_04369_),
    .ZN(_06071_));
 NOR2_X1 _23093_ (.A1(_04391_),
    .A2(_06071_),
    .ZN(_06072_));
 NAND2_X1 _23094_ (.A1(_04308_),
    .A2(_05119_),
    .ZN(_06073_));
 NAND2_X1 _23095_ (.A1(_04723_),
    .A2(_05867_),
    .ZN(_06074_));
 AOI21_X2 _23096_ (.A(_04342_),
    .B1(_06073_),
    .B2(_06074_),
    .ZN(_06075_));
 AND2_X1 _23097_ (.A1(_15565_),
    .A2(_05079_),
    .ZN(_06076_));
 INV_X1 _23098_ (.A(_15738_),
    .ZN(_06077_));
 NAND2_X4 _23099_ (.A1(_04498_),
    .A2(_06077_),
    .ZN(_06078_));
 AND2_X4 _23100_ (.A1(_15745_),
    .A2(_06078_),
    .ZN(_06079_));
 NOR2_X1 _23101_ (.A1(_15745_),
    .A2(_06078_),
    .ZN(_06080_));
 NOR3_X2 _23102_ (.A1(_05079_),
    .A2(_06079_),
    .A3(_06080_),
    .ZN(_06081_));
 NOR3_X4 _23103_ (.A1(_04622_),
    .A2(_06076_),
    .A3(_06081_),
    .ZN(_06082_));
 AND2_X1 _23104_ (.A1(_04622_),
    .A2(_03804_),
    .ZN(_06083_));
 NOR3_X4 _23105_ (.A1(_11408_),
    .A2(_06082_),
    .A3(_06083_),
    .ZN(_06084_));
 AOI222_X2 _23106_ (.A1(net143),
    .A2(_04518_),
    .B1(_05074_),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .C1(\cs_registers_i.mscratch_q[18] ),
    .C2(_04523_),
    .ZN(_06085_));
 AOI22_X1 _23107_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(_04771_),
    .B1(_04514_),
    .B2(\cs_registers_i.mie_q[2] ),
    .ZN(_06086_));
 AOI22_X1 _23108_ (.A1(net80),
    .A2(_04528_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .ZN(_06087_));
 OAI21_X1 _23109_ (.A(_04533_),
    .B1(_04536_),
    .B2(_01175_),
    .ZN(_06088_));
 AOI221_X1 _23110_ (.A(_06088_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[18] ),
    .C1(\cs_registers_i.dscratch1_q[18] ),
    .C2(_04529_),
    .ZN(_06089_));
 AND4_X1 _23111_ (.A1(_06085_),
    .A2(_06086_),
    .A3(_06087_),
    .A4(_06089_),
    .ZN(_06090_));
 BUF_X2 _23112_ (.A(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .Z(_06091_));
 BUF_X2 _23113_ (.A(\cs_registers_i.mhpmcounter[2][50] ),
    .Z(_06092_));
 AOI22_X2 _23114_ (.A1(_06091_),
    .A2(_04963_),
    .B1(_04964_),
    .B2(_06092_),
    .ZN(_06093_));
 BUF_X2 _23115_ (.A(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .Z(_06094_));
 CLKBUF_X2 _23116_ (.A(\cs_registers_i.mhpmcounter[2][18] ),
    .Z(_06095_));
 AOI22_X2 _23117_ (.A1(_06094_),
    .A2(_04963_),
    .B1(_04964_),
    .B2(_06095_),
    .ZN(_06096_));
 OAI221_X2 _23118_ (.A(_06090_),
    .B1(_06093_),
    .B2(_05031_),
    .C1(_04560_),
    .C2(_06096_),
    .ZN(_06097_));
 NOR4_X4 _23119_ (.A1(_06072_),
    .A2(_06075_),
    .A3(_06084_),
    .A4(_06097_),
    .ZN(_06098_));
 AOI21_X4 _23120_ (.A(_06067_),
    .B1(_06098_),
    .B2(_04764_),
    .ZN(_06099_));
 BUF_X2 _23121_ (.A(_06099_),
    .Z(_06100_));
 MUX2_X1 _23122_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .S(_05929_),
    .Z(_01216_));
 NAND2_X1 _23123_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .A2(_05416_),
    .ZN(_06101_));
 OR2_X1 _23124_ (.A1(_05949_),
    .A2(_05828_),
    .ZN(_06102_));
 AOI221_X1 _23125_ (.A(_04352_),
    .B1(_04360_),
    .B2(_15991_),
    .C1(_04363_),
    .C2(_15990_),
    .ZN(_06103_));
 AOI21_X1 _23126_ (.A(_06103_),
    .B1(_04370_),
    .B2(_15994_),
    .ZN(_06104_));
 AOI21_X2 _23127_ (.A(_06104_),
    .B1(_04825_),
    .B2(\alu_adder_result_ex[19] ),
    .ZN(_06105_));
 INV_X1 _23128_ (.A(_15580_),
    .ZN(_06106_));
 OAI21_X2 _23129_ (.A(_12102_),
    .B1(_06106_),
    .B2(_04502_),
    .ZN(_06107_));
 NAND2_X1 _23130_ (.A1(_04472_),
    .A2(_06025_),
    .ZN(_06108_));
 AOI21_X2 _23131_ (.A(_04466_),
    .B1(_04636_),
    .B2(_06108_),
    .ZN(_06109_));
 XOR2_X2 _23132_ (.A(_15751_),
    .B(_06109_),
    .Z(_06110_));
 AOI21_X4 _23133_ (.A(_06107_),
    .B1(_06110_),
    .B2(_04791_),
    .ZN(_06111_));
 OAI21_X2 _23134_ (.A(_03449_),
    .B1(_03806_),
    .B2(_12103_),
    .ZN(_06112_));
 OAI22_X4 _23135_ (.A1(_04391_),
    .A2(_06105_),
    .B1(_06111_),
    .B2(_06112_),
    .ZN(_06113_));
 NOR2_X1 _23136_ (.A1(_01176_),
    .A2(_04728_),
    .ZN(_06114_));
 AOI221_X2 _23137_ (.A(_06114_),
    .B1(_04731_),
    .B2(\cs_registers_i.dscratch0_q[19] ),
    .C1(\cs_registers_i.mie_q[3] ),
    .C2(_04733_),
    .ZN(_06115_));
 AOI22_X2 _23138_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_04736_),
    .B1(_04738_),
    .B2(\cs_registers_i.mscratch_q[19] ),
    .ZN(_06116_));
 AOI221_X2 _23139_ (.A(_04741_),
    .B1(_04742_),
    .B2(net144),
    .C1(net81),
    .C2(_04743_),
    .ZN(_06117_));
 NAND3_X2 _23140_ (.A1(_06115_),
    .A2(_06116_),
    .A3(_06117_),
    .ZN(_06118_));
 AOI222_X2 _23141_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_04747_),
    .B1(_04748_),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .C1(_04749_),
    .C2(\cs_registers_i.dscratch1_q[19] ),
    .ZN(_06119_));
 BUF_X2 _23142_ (.A(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .Z(_06120_));
 AOI22_X2 _23143_ (.A1(_06120_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(\cs_registers_i.mhpmcounter[2][51] ),
    .ZN(_06121_));
 OAI21_X1 _23144_ (.A(_06119_),
    .B1(_06121_),
    .B2(_04756_),
    .ZN(_06122_));
 BUF_X2 _23145_ (.A(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .Z(_06123_));
 CLKBUF_X2 _23146_ (.A(\cs_registers_i.mhpmcounter[2][19] ),
    .Z(_06124_));
 AOI22_X2 _23147_ (.A1(_06123_),
    .A2(_04550_),
    .B1(_04553_),
    .B2(_06124_),
    .ZN(_06125_));
 NOR2_X1 _23148_ (.A1(_03532_),
    .A2(_06125_),
    .ZN(_06126_));
 OR3_X4 _23149_ (.A1(_06118_),
    .A2(_06122_),
    .A3(_06126_),
    .ZN(_06127_));
 NOR3_X4 _23150_ (.A1(_04342_),
    .A2(_04723_),
    .A3(_05830_),
    .ZN(_06128_));
 NOR3_X4 _23151_ (.A1(_06113_),
    .A2(_06127_),
    .A3(_06128_),
    .ZN(_06129_));
 OAI21_X1 _23152_ (.A(_05982_),
    .B1(_05055_),
    .B2(_04308_),
    .ZN(_06130_));
 NAND2_X1 _23153_ (.A1(_04276_),
    .A2(_06130_),
    .ZN(_06131_));
 NAND4_X4 _23154_ (.A1(_04600_),
    .A2(_06102_),
    .A3(_06129_),
    .A4(_06131_),
    .ZN(_06132_));
 NAND3_X1 _23155_ (.A1(_05421_),
    .A2(_05503_),
    .A3(_05507_),
    .ZN(_06133_));
 MUX2_X1 _23156_ (.A(net48),
    .B(\load_store_unit_i.rdata_q[27] ),
    .S(_04594_),
    .Z(_06134_));
 OAI21_X1 _23157_ (.A(_06133_),
    .B1(_06134_),
    .B2(_04597_),
    .ZN(_06135_));
 OAI21_X1 _23158_ (.A(_04616_),
    .B1(_04859_),
    .B2(_06135_),
    .ZN(_06136_));
 OAI21_X2 _23159_ (.A(_06132_),
    .B1(_06136_),
    .B2(_04764_),
    .ZN(_06137_));
 CLKBUF_X3 _23160_ (.A(_06137_),
    .Z(_06138_));
 OAI21_X1 _23161_ (.A(_06101_),
    .B1(_06138_),
    .B2(_05465_),
    .ZN(_01217_));
 NAND3_X1 _23162_ (.A1(_04596_),
    .A2(_05515_),
    .A3(_05519_),
    .ZN(_06139_));
 MUX2_X1 _23163_ (.A(net50),
    .B(\load_store_unit_i.rdata_q[28] ),
    .S(_04586_),
    .Z(_06140_));
 OAI21_X1 _23164_ (.A(_06139_),
    .B1(_06140_),
    .B2(_05421_),
    .ZN(_06141_));
 INV_X1 _23165_ (.A(_06141_),
    .ZN(_06142_));
 AOI21_X4 _23166_ (.A(_04617_),
    .B1(_06142_),
    .B2(_04583_),
    .ZN(_06143_));
 NOR2_X1 _23167_ (.A1(_15998_),
    .A2(_04664_),
    .ZN(_06144_));
 MUX2_X1 _23168_ (.A(_15999_),
    .B(_16002_),
    .S(_04362_),
    .Z(_06145_));
 AOI21_X1 _23169_ (.A(_06144_),
    .B1(_06145_),
    .B2(_04664_),
    .ZN(_06146_));
 OAI21_X1 _23170_ (.A(_05116_),
    .B1(_06146_),
    .B2(_04387_),
    .ZN(_06147_));
 AOI221_X1 _23171_ (.A(_06147_),
    .B1(_05120_),
    .B2(_04831_),
    .C1(\alu_adder_result_ex[20] ),
    .C2(_04369_),
    .ZN(_06148_));
 NOR2_X1 _23172_ (.A1(_04391_),
    .A2(_06148_),
    .ZN(_06149_));
 AOI21_X1 _23173_ (.A(_11407_),
    .B1(_03808_),
    .B2(_04622_),
    .ZN(_06150_));
 OAI21_X4 _23174_ (.A(_15751_),
    .B1(_06079_),
    .B2(_15744_),
    .ZN(_06151_));
 NAND2_X2 _23175_ (.A1(_06151_),
    .A2(_04635_),
    .ZN(_06152_));
 XNOR2_X2 _23176_ (.A(_06152_),
    .B(_04465_),
    .ZN(_06153_));
 MUX2_X1 _23177_ (.A(_15588_),
    .B(_06153_),
    .S(_04502_),
    .Z(_06154_));
 OAI21_X4 _23178_ (.A(_06150_),
    .B1(net304),
    .B2(_06154_),
    .ZN(_06155_));
 INV_X4 _23179_ (.A(_06155_),
    .ZN(_06156_));
 AOI22_X1 _23180_ (.A1(\cs_registers_i.mscratch_q[20] ),
    .A2(_04524_),
    .B1(_04521_),
    .B2(\cs_registers_i.mtval_q[20] ),
    .ZN(_06157_));
 AOI22_X1 _23181_ (.A1(net145),
    .A2(_04518_),
    .B1(_04544_),
    .B2(\cs_registers_i.csr_mepc_o[20] ),
    .ZN(_06158_));
 NAND2_X1 _23182_ (.A1(_06157_),
    .A2(_06158_),
    .ZN(_06159_));
 AOI22_X1 _23183_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(_04515_),
    .B1(_04530_),
    .B2(\cs_registers_i.dscratch1_q[20] ),
    .ZN(_06160_));
 AOI22_X1 _23184_ (.A1(net83),
    .A2(_04528_),
    .B1(_04968_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .ZN(_06161_));
 NAND2_X1 _23185_ (.A1(_06160_),
    .A2(_06161_),
    .ZN(_06162_));
 NAND2_X1 _23186_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_04511_),
    .ZN(_06163_));
 OR2_X1 _23187_ (.A1(_01177_),
    .A2(_04537_),
    .ZN(_06164_));
 NAND3_X1 _23188_ (.A1(_04247_),
    .A2(_06163_),
    .A3(_06164_),
    .ZN(_06165_));
 NOR3_X2 _23189_ (.A1(_06159_),
    .A2(_06162_),
    .A3(_06165_),
    .ZN(_06166_));
 AOI22_X2 _23190_ (.A1(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .A2(_04959_),
    .B1(_04960_),
    .B2(\cs_registers_i.mhpmcounter[2][52] ),
    .ZN(_06167_));
 BUF_X2 _23191_ (.A(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .Z(_06168_));
 AOI22_X2 _23192_ (.A1(_06168_),
    .A2(_04551_),
    .B1(_04554_),
    .B2(\cs_registers_i.mhpmcounter[2][20] ),
    .ZN(_06169_));
 OAI221_X2 _23193_ (.A(_06166_),
    .B1(_06167_),
    .B2(_05031_),
    .C1(_04560_),
    .C2(_06169_),
    .ZN(_06170_));
 NOR3_X2 _23194_ (.A1(_04725_),
    .A2(_05796_),
    .A3(_05798_),
    .ZN(_06171_));
 NOR4_X4 _23195_ (.A1(_06149_),
    .A2(_06156_),
    .A3(_06170_),
    .A4(_06171_),
    .ZN(_06172_));
 AOI21_X4 _23196_ (.A(_06143_),
    .B1(_04600_),
    .B2(_06172_),
    .ZN(_06173_));
 BUF_X4 _23197_ (.A(_06173_),
    .Z(_06174_));
 MUX2_X1 _23198_ (.A(_06174_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .S(_05929_),
    .Z(_01218_));
 NAND3_X1 _23199_ (.A1(_04596_),
    .A2(_05548_),
    .A3(_05552_),
    .ZN(_06175_));
 MUX2_X1 _23200_ (.A(net51),
    .B(\load_store_unit_i.rdata_q[29] ),
    .S(_04586_),
    .Z(_06176_));
 OAI21_X1 _23201_ (.A(_06175_),
    .B1(_06176_),
    .B2(_05421_),
    .ZN(_06177_));
 INV_X1 _23202_ (.A(_06177_),
    .ZN(_06178_));
 AOI21_X4 _23203_ (.A(_04617_),
    .B1(_06178_),
    .B2(_04582_),
    .ZN(_06179_));
 NAND3_X1 _23204_ (.A1(_04633_),
    .A2(_04634_),
    .A3(_04654_),
    .ZN(_06180_));
 NOR2_X1 _23205_ (.A1(_04625_),
    .A2(_04655_),
    .ZN(_06181_));
 NAND2_X1 _23206_ (.A1(_06180_),
    .A2(_06181_),
    .ZN(_06182_));
 AOI21_X2 _23207_ (.A(net304),
    .B1(_14126_),
    .B2(_05079_),
    .ZN(_06183_));
 AOI221_X2 _23208_ (.A(_11407_),
    .B1(_06182_),
    .B2(_06183_),
    .C1(_00845_),
    .C2(_04622_),
    .ZN(_06184_));
 AOI22_X1 _23209_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(_04523_),
    .B1(_04543_),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .ZN(_06185_));
 AOI22_X1 _23210_ (.A1(net146),
    .A2(_04517_),
    .B1(_04520_),
    .B2(\cs_registers_i.mtval_q[21] ),
    .ZN(_06186_));
 AND2_X1 _23211_ (.A1(_06185_),
    .A2(_06186_),
    .ZN(_06187_));
 AOI222_X2 _23212_ (.A1(\cs_registers_i.dscratch0_q[21] ),
    .A2(_04771_),
    .B1(_04775_),
    .B2(\cs_registers_i.dscratch1_q[21] ),
    .C1(\cs_registers_i.csr_mstatus_tw_o ),
    .C2(_05487_),
    .ZN(_06188_));
 OAI21_X1 _23213_ (.A(_04534_),
    .B1(_04537_),
    .B2(_01178_),
    .ZN(_06189_));
 AOI21_X1 _23214_ (.A(_06189_),
    .B1(_04515_),
    .B2(\cs_registers_i.mie_q[5] ),
    .ZN(_06190_));
 AOI22_X1 _23215_ (.A1(net84),
    .A2(_04528_),
    .B1(_04773_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .ZN(_06191_));
 AND4_X1 _23216_ (.A1(_06187_),
    .A2(_06188_),
    .A3(_06190_),
    .A4(_06191_),
    .ZN(_06192_));
 BUF_X2 _23217_ (.A(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .Z(_06193_));
 BUF_X2 _23218_ (.A(\cs_registers_i.mhpmcounter[2][53] ),
    .Z(_06194_));
 AOI22_X4 _23219_ (.A1(_06193_),
    .A2(_04784_),
    .B1(_04785_),
    .B2(_06194_),
    .ZN(_06195_));
 AOI22_X2 _23220_ (.A1(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\cs_registers_i.mhpmcounter[2][21] ),
    .ZN(_06196_));
 OAI221_X2 _23221_ (.A(_06192_),
    .B1(_06195_),
    .B2(_04557_),
    .C1(_04783_),
    .C2(_06196_),
    .ZN(_06197_));
 INV_X1 _23222_ (.A(_16006_),
    .ZN(_06198_));
 AOI22_X1 _23223_ (.A1(_06198_),
    .A2(_04352_),
    .B1(_04368_),
    .B2(\alu_adder_result_ex[21] ),
    .ZN(_06199_));
 AOI22_X1 _23224_ (.A1(_16007_),
    .A2(_04360_),
    .B1(_04983_),
    .B2(_16010_),
    .ZN(_06200_));
 OAI21_X1 _23225_ (.A(_06199_),
    .B1(_06200_),
    .B2(_04353_),
    .ZN(_06201_));
 AOI221_X1 _23226_ (.A(_06201_),
    .B1(_05120_),
    .B2(_05009_),
    .C1(_04307_),
    .C2(_05868_),
    .ZN(_06202_));
 NOR2_X1 _23227_ (.A1(_04391_),
    .A2(_06202_),
    .ZN(_06203_));
 AND3_X1 _23228_ (.A1(_04457_),
    .A2(_04459_),
    .A3(_05733_),
    .ZN(_06204_));
 NOR4_X4 _23229_ (.A1(_06184_),
    .A2(_06197_),
    .A3(_06203_),
    .A4(_06204_),
    .ZN(_06205_));
 AOI21_X4 _23230_ (.A(_06179_),
    .B1(_06205_),
    .B2(_04600_),
    .ZN(_06206_));
 BUF_X2 _23231_ (.A(_06206_),
    .Z(_06207_));
 MUX2_X1 _23232_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .S(_05929_),
    .Z(_01219_));
 BUF_X4 _23233_ (.A(_05210_),
    .Z(_06208_));
 MUX2_X1 _23234_ (.A(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .B(_06208_),
    .S(_05415_),
    .Z(_01220_));
 MUX2_X1 _23235_ (.A(_04602_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .S(_05929_),
    .Z(_01221_));
 MUX2_X1 _23236_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .S(_05929_),
    .Z(_01222_));
 NAND2_X1 _23237_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .A2(_05416_),
    .ZN(_06209_));
 OAI21_X1 _23238_ (.A(_06209_),
    .B1(_05465_),
    .B2(_04908_),
    .ZN(_01223_));
 NAND2_X1 _23239_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .A2(_05416_),
    .ZN(_06210_));
 OAI21_X4 _23240_ (.A(_06210_),
    .B1(net442),
    .B2(_05465_),
    .ZN(_01224_));
 MUX2_X1 _23241_ (.A(net418),
    .B(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .S(_05929_),
    .Z(_01225_));
 MUX2_X1 _23242_ (.A(net333),
    .B(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .S(_05929_),
    .Z(_01226_));
 MUX2_X1 _23243_ (.A(net409),
    .B(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .S(_05375_),
    .Z(_01227_));
 NAND2_X1 _23244_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A2(_05416_),
    .ZN(_06211_));
 OAI21_X4 _23245_ (.A(_06211_),
    .B1(net445),
    .B2(_05465_),
    .ZN(_01228_));
 MUX2_X1 _23246_ (.A(_05211_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .S(_05375_),
    .Z(_01229_));
 NAND2_X1 _23247_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A2(_05416_),
    .ZN(_06212_));
 OAI21_X2 _23248_ (.A(_06212_),
    .B1(net441),
    .B2(_05465_),
    .ZN(_01230_));
 NAND2_X1 _23249_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .A2(_05803_),
    .ZN(_06213_));
 OAI21_X4 _23250_ (.A(_06213_),
    .B1(net441),
    .B2(_05806_),
    .ZN(_01231_));
 NOR2_X4 _23251_ (.A1(_04603_),
    .A2(_04851_),
    .ZN(_06214_));
 NAND2_X4 _23252_ (.A1(_04613_),
    .A2(_06214_),
    .ZN(_06215_));
 BUF_X8 _23253_ (.A(_06215_),
    .Z(_06216_));
 MUX2_X1 _23254_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(_06216_),
    .Z(_01232_));
 MUX2_X1 _23255_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S(_06216_),
    .Z(_01233_));
 BUF_X4 _23256_ (.A(_06215_),
    .Z(_06217_));
 NAND2_X1 _23257_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .A2(_06217_),
    .ZN(_06218_));
 BUF_X4 _23258_ (.A(_06215_),
    .Z(_06219_));
 OAI21_X1 _23259_ (.A(_06218_),
    .B1(_06219_),
    .B2(_05464_),
    .ZN(_01234_));
 NAND2_X1 _23260_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .A2(_06217_),
    .ZN(_06220_));
 OAI21_X1 _23261_ (.A(_06220_),
    .B1(_06219_),
    .B2(_05510_),
    .ZN(_01235_));
 MUX2_X1 _23262_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S(_06216_),
    .Z(_01236_));
 MUX2_X1 _23263_ (.A(_05580_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S(_06216_),
    .Z(_01237_));
 MUX2_X1 _23264_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S(_06216_),
    .Z(_01238_));
 MUX2_X1 _23265_ (.A(_05653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S(_06216_),
    .Z(_01239_));
 NAND2_X1 _23266_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .A2(_06217_),
    .ZN(_06221_));
 BUF_X4 _23267_ (.A(_05687_),
    .Z(_06222_));
 OAI21_X1 _23268_ (.A(_06221_),
    .B1(_06219_),
    .B2(_06222_),
    .ZN(_01240_));
 MUX2_X1 _23269_ (.A(_05721_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S(_06216_),
    .Z(_01241_));
 BUF_X2 _23270_ (.A(_05371_),
    .Z(_06223_));
 BUF_X8 _23271_ (.A(_05412_),
    .Z(_06224_));
 AOI21_X4 _23272_ (.A(_10899_),
    .B1(_04605_),
    .B2(_04611_),
    .ZN(_06225_));
 BUF_X8 _23273_ (.A(_06225_),
    .Z(_06226_));
 AND3_X1 _23274_ (.A1(_06224_),
    .A2(_10904_),
    .A3(_06226_),
    .ZN(_06227_));
 BUF_X4 _23275_ (.A(_06227_),
    .Z(_06228_));
 BUF_X4 _23276_ (.A(_06228_),
    .Z(_06229_));
 MUX2_X1 _23277_ (.A(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .B(_06223_),
    .S(_06229_),
    .Z(_01242_));
 MUX2_X1 _23278_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S(_06216_),
    .Z(_01243_));
 MUX2_X1 _23279_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S(_06216_),
    .Z(_01244_));
 NAND2_X1 _23280_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .A2(_06217_),
    .ZN(_06230_));
 CLKBUF_X3 _23281_ (.A(_05849_),
    .Z(_06231_));
 OAI21_X1 _23282_ (.A(_06230_),
    .B1(_06219_),
    .B2(_06231_),
    .ZN(_01245_));
 MUX2_X1 _23283_ (.A(_05890_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S(_06216_),
    .Z(_01246_));
 BUF_X4 _23284_ (.A(_06215_),
    .Z(_06232_));
 MUX2_X1 _23285_ (.A(_05928_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S(_06232_),
    .Z(_01247_));
 MUX2_X1 _23286_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S(_06232_),
    .Z(_01248_));
 NAND2_X1 _23287_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .A2(_06217_),
    .ZN(_06233_));
 CLKBUF_X3 _23288_ (.A(_06015_),
    .Z(_06234_));
 OAI21_X1 _23289_ (.A(_06233_),
    .B1(_06219_),
    .B2(_06234_),
    .ZN(_01249_));
 MUX2_X1 _23290_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S(_06232_),
    .Z(_01250_));
 MUX2_X1 _23291_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S(_06232_),
    .Z(_01251_));
 NAND2_X1 _23292_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .A2(_06217_),
    .ZN(_06235_));
 OAI21_X1 _23293_ (.A(_06235_),
    .B1(_06219_),
    .B2(_06138_),
    .ZN(_01252_));
 BUF_X2 _23294_ (.A(_05409_),
    .Z(_06236_));
 MUX2_X1 _23295_ (.A(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .B(_06236_),
    .S(_06229_),
    .Z(_01253_));
 MUX2_X1 _23296_ (.A(net405),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S(_06232_),
    .Z(_01254_));
 MUX2_X1 _23297_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S(_06232_),
    .Z(_01255_));
 MUX2_X1 _23298_ (.A(_04602_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S(_06232_),
    .Z(_01256_));
 MUX2_X1 _23299_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S(_06232_),
    .Z(_01257_));
 NAND2_X1 _23300_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .A2(_06217_),
    .ZN(_06237_));
 OAI21_X1 _23301_ (.A(_06237_),
    .B1(_06219_),
    .B2(_04908_),
    .ZN(_01258_));
 NAND2_X1 _23302_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .A2(_06217_),
    .ZN(_06238_));
 OAI21_X4 _23303_ (.A(_06238_),
    .B1(net442),
    .B2(_06219_),
    .ZN(_01259_));
 MUX2_X1 _23304_ (.A(net418),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S(_06232_),
    .Z(_01260_));
 MUX2_X1 _23305_ (.A(_04850_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S(_06232_),
    .Z(_01261_));
 MUX2_X1 _23306_ (.A(net409),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S(_06215_),
    .Z(_01262_));
 NAND2_X1 _23307_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .A2(_06217_),
    .ZN(_06239_));
 OAI21_X4 _23308_ (.A(_06239_),
    .B1(net445),
    .B2(_06219_),
    .ZN(_01263_));
 NAND3_X4 _23309_ (.A1(_06224_),
    .A2(_10904_),
    .A3(_06226_),
    .ZN(_06240_));
 BUF_X4 _23310_ (.A(_06240_),
    .Z(_06241_));
 NAND2_X1 _23311_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .A2(_06241_),
    .ZN(_06242_));
 OAI21_X1 _23312_ (.A(_06242_),
    .B1(_06241_),
    .B2(_05464_),
    .ZN(_01264_));
 MUX2_X1 _23313_ (.A(net400),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S(_06215_),
    .Z(_01265_));
 NAND2_X1 _23314_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .A2(_06217_),
    .ZN(_06243_));
 OAI21_X4 _23315_ (.A(_06243_),
    .B1(net441),
    .B2(_06219_),
    .ZN(_01266_));
 NAND2_X1 _23316_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .A2(_06241_),
    .ZN(_06244_));
 OAI21_X1 _23317_ (.A(_06244_),
    .B1(_06241_),
    .B2(_05510_),
    .ZN(_01267_));
 NOR3_X4 _23318_ (.A1(_10394_),
    .A2(_11315_),
    .A3(_10903_),
    .ZN(_06245_));
 NAND2_X4 _23319_ (.A1(_04854_),
    .A2(_06245_),
    .ZN(_06246_));
 MUX2_X1 _23320_ (.A(_05721_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .S(_06246_),
    .Z(_01268_));
 NAND2_X1 _23321_ (.A1(_05314_),
    .A2(_05316_),
    .ZN(_06247_));
 NOR4_X4 _23322_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_03627_),
    .A3(_03637_),
    .A4(_03642_),
    .ZN(_06248_));
 NOR4_X4 _23323_ (.A1(\alu_adder_result_ex[22] ),
    .A2(\alu_adder_result_ex[24] ),
    .A3(\alu_adder_result_ex[31] ),
    .A4(_03644_),
    .ZN(_06249_));
 NAND3_X2 _23324_ (.A1(_06248_),
    .A2(_06249_),
    .A3(_05314_),
    .ZN(_06250_));
 NAND3_X4 _23325_ (.A1(_10350_),
    .A2(_10909_),
    .A3(_11427_),
    .ZN(_06251_));
 NOR3_X4 _23326_ (.A1(net307),
    .A2(_03434_),
    .A3(_06251_),
    .ZN(_06252_));
 NAND3_X4 _23327_ (.A1(_06247_),
    .A2(_06250_),
    .A3(_06252_),
    .ZN(_06253_));
 NOR2_X1 _23328_ (.A1(_10305_),
    .A2(_10909_),
    .ZN(_06254_));
 OAI21_X1 _23329_ (.A(_06254_),
    .B1(_03456_),
    .B2(_10350_),
    .ZN(_06255_));
 NOR2_X2 _23330_ (.A1(_10909_),
    .A2(_03434_),
    .ZN(_06256_));
 AOI21_X2 _23331_ (.A(_04229_),
    .B1(_06256_),
    .B2(_03456_),
    .ZN(_06257_));
 NOR2_X1 _23332_ (.A1(_10350_),
    .A2(_03438_),
    .ZN(_06258_));
 OAI21_X1 _23333_ (.A(_10332_),
    .B1(_10340_),
    .B2(_03884_),
    .ZN(_06259_));
 OAI21_X1 _23334_ (.A(_06258_),
    .B1(_06259_),
    .B2(_11401_),
    .ZN(_06260_));
 NOR2_X1 _23335_ (.A1(_03885_),
    .A2(_04229_),
    .ZN(_06261_));
 OAI221_X2 _23336_ (.A(_06255_),
    .B1(_06257_),
    .B2(_06260_),
    .C1(_06261_),
    .C2(_06251_),
    .ZN(_06262_));
 NOR3_X4 _23337_ (.A1(_03643_),
    .A2(_03645_),
    .A3(_05327_),
    .ZN(_06263_));
 AOI22_X4 _23338_ (.A1(_11418_),
    .A2(_06262_),
    .B1(_06252_),
    .B2(_06263_),
    .ZN(_06264_));
 NAND2_X4 _23339_ (.A1(_06253_),
    .A2(_06264_),
    .ZN(_06265_));
 AND2_X1 _23340_ (.A1(_03869_),
    .A2(_03872_),
    .ZN(_06266_));
 AOI21_X1 _23341_ (.A(net69),
    .B1(_03879_),
    .B2(_10304_),
    .ZN(_06267_));
 OR2_X2 _23342_ (.A1(_03954_),
    .A2(_06267_),
    .ZN(_06268_));
 NAND3_X1 _23343_ (.A1(_03458_),
    .A2(_11423_),
    .A3(_06268_),
    .ZN(_06269_));
 NOR3_X1 _23344_ (.A1(_11420_),
    .A2(_06266_),
    .A3(_06269_),
    .ZN(_06270_));
 NAND2_X1 _23345_ (.A1(_03894_),
    .A2(_03895_),
    .ZN(_06271_));
 OR2_X1 _23346_ (.A1(\id_stage_i.controller_i.load_err_d ),
    .A2(\id_stage_i.controller_i.store_err_d ),
    .ZN(_06272_));
 NOR4_X1 _23347_ (.A1(_10468_),
    .A2(_15525_),
    .A3(_10876_),
    .A4(_10980_),
    .ZN(_06273_));
 INV_X1 _23348_ (.A(_15525_),
    .ZN(_06274_));
 NOR3_X1 _23349_ (.A1(_15527_),
    .A2(_06274_),
    .A3(_10891_),
    .ZN(_06275_));
 AOI21_X1 _23350_ (.A(_06273_),
    .B1(_06275_),
    .B2(_03475_),
    .ZN(_06276_));
 NOR3_X1 _23351_ (.A1(_10885_),
    .A2(_03486_),
    .A3(_06276_),
    .ZN(_06277_));
 NOR4_X1 _23352_ (.A1(_03472_),
    .A2(_06271_),
    .A3(_06272_),
    .A4(_06277_),
    .ZN(_06278_));
 AND3_X1 _23353_ (.A1(_03479_),
    .A2(_03610_),
    .A3(_06278_),
    .ZN(_06279_));
 OAI211_X2 _23354_ (.A(_03509_),
    .B(_06279_),
    .C1(_03603_),
    .C2(_03552_),
    .ZN(_06280_));
 AND3_X1 _23355_ (.A1(_01161_),
    .A2(_03479_),
    .A3(_03610_),
    .ZN(_06281_));
 OAI21_X1 _23356_ (.A(_06278_),
    .B1(_06281_),
    .B2(_03461_),
    .ZN(_06282_));
 AND2_X1 _23357_ (.A1(_06280_),
    .A2(_06282_),
    .ZN(_06283_));
 NOR2_X1 _23358_ (.A1(_11426_),
    .A2(_06283_),
    .ZN(_06284_));
 OAI21_X1 _23359_ (.A(_06284_),
    .B1(_06268_),
    .B2(_06265_),
    .ZN(_06285_));
 NOR3_X2 _23360_ (.A1(_03477_),
    .A2(_03869_),
    .A3(_03880_),
    .ZN(_06286_));
 NAND3_X2 _23361_ (.A1(_11421_),
    .A2(_03875_),
    .A3(_11424_),
    .ZN(_06287_));
 NOR2_X1 _23362_ (.A1(_03436_),
    .A2(_06287_),
    .ZN(_06288_));
 AND2_X1 _23363_ (.A1(_06286_),
    .A2(_06288_),
    .ZN(_06289_));
 NOR2_X1 _23364_ (.A1(_03954_),
    .A2(_06267_),
    .ZN(_06290_));
 NAND3_X2 _23365_ (.A1(_11933_),
    .A2(_03609_),
    .A3(_03851_),
    .ZN(_06291_));
 NOR2_X1 _23366_ (.A1(_03848_),
    .A2(_03847_),
    .ZN(_06292_));
 AOI21_X2 _23367_ (.A(_06292_),
    .B1(_03464_),
    .B2(\cs_registers_i.dcsr_q[15] ),
    .ZN(_06293_));
 OAI21_X1 _23368_ (.A(_06290_),
    .B1(_06291_),
    .B2(_06293_),
    .ZN(_06294_));
 NAND2_X1 _23369_ (.A1(_03461_),
    .A2(_06294_),
    .ZN(_06295_));
 NOR2_X1 _23370_ (.A1(_03891_),
    .A2(_06271_),
    .ZN(_06296_));
 AOI21_X2 _23371_ (.A(_06295_),
    .B1(_06296_),
    .B2(_03472_),
    .ZN(_06297_));
 NOR3_X1 _23372_ (.A1(_03436_),
    .A2(_03458_),
    .A3(_11424_),
    .ZN(_06298_));
 OAI21_X1 _23373_ (.A(_11423_),
    .B1(_06290_),
    .B2(_11421_),
    .ZN(_06299_));
 AOI21_X1 _23374_ (.A(_06298_),
    .B1(_06299_),
    .B2(_03436_),
    .ZN(_06300_));
 OAI21_X1 _23375_ (.A(_03890_),
    .B1(_06300_),
    .B2(_11422_),
    .ZN(_06301_));
 NOR3_X1 _23376_ (.A1(_06289_),
    .A2(_06297_),
    .A3(_06301_),
    .ZN(_06302_));
 AOI222_X2 _23377_ (.A1(_11422_),
    .A2(_03877_),
    .B1(_06265_),
    .B2(_06270_),
    .C1(_06285_),
    .C2(_06302_),
    .ZN(_01269_));
 NAND2_X1 _23378_ (.A1(_03869_),
    .A2(_03872_),
    .ZN(_06303_));
 NOR2_X1 _23379_ (.A1(_06265_),
    .A2(_06303_),
    .ZN(_06304_));
 OAI221_X1 _23380_ (.A(_03931_),
    .B1(_06265_),
    .B2(_06268_),
    .C1(_06304_),
    .C2(_11421_),
    .ZN(_06305_));
 NAND3_X2 _23381_ (.A1(_03931_),
    .A2(_06280_),
    .A3(_06282_),
    .ZN(_06306_));
 NOR2_X1 _23382_ (.A1(_03840_),
    .A2(_06295_),
    .ZN(_06307_));
 NAND3_X1 _23383_ (.A1(_10304_),
    .A2(_06266_),
    .A3(_06277_),
    .ZN(_06308_));
 NAND3_X1 _23384_ (.A1(_03605_),
    .A2(_10678_),
    .A3(_10882_),
    .ZN(_06309_));
 OAI21_X1 _23385_ (.A(_06308_),
    .B1(_06309_),
    .B2(_03465_),
    .ZN(_06310_));
 OAI22_X1 _23386_ (.A1(_03458_),
    .A2(_11423_),
    .B1(_06303_),
    .B2(_06269_),
    .ZN(_06311_));
 AOI221_X2 _23387_ (.A(_06289_),
    .B1(_06307_),
    .B2(_06310_),
    .C1(_06311_),
    .C2(_04160_),
    .ZN(_06312_));
 NAND3_X1 _23388_ (.A1(_06305_),
    .A2(_06306_),
    .A3(_06312_),
    .ZN(_01270_));
 NAND3_X1 _23389_ (.A1(_11423_),
    .A2(_04160_),
    .A3(_06268_),
    .ZN(_06313_));
 OAI21_X1 _23390_ (.A(_06313_),
    .B1(_11423_),
    .B2(_03875_),
    .ZN(_06314_));
 NAND2_X1 _23391_ (.A1(_11421_),
    .A2(_03875_),
    .ZN(_06315_));
 NAND2_X1 _23392_ (.A1(_06315_),
    .A2(_03877_),
    .ZN(_06316_));
 AOI222_X2 _23393_ (.A1(_03854_),
    .A2(_06297_),
    .B1(_06314_),
    .B2(_03458_),
    .C1(_11420_),
    .C2(_06316_),
    .ZN(_06317_));
 OR2_X1 _23394_ (.A1(_06265_),
    .A2(_06283_),
    .ZN(_06318_));
 OAI21_X1 _23395_ (.A(_03931_),
    .B1(_06268_),
    .B2(_06318_),
    .ZN(_06319_));
 AOI221_X1 _23396_ (.A(_06289_),
    .B1(_06317_),
    .B2(_06319_),
    .C1(_03877_),
    .C2(_11422_),
    .ZN(_01271_));
 NAND2_X1 _23397_ (.A1(_11425_),
    .A2(_06290_),
    .ZN(_06320_));
 AOI21_X1 _23398_ (.A(_06320_),
    .B1(_06318_),
    .B2(_11420_),
    .ZN(_06321_));
 AOI21_X1 _23399_ (.A(_03952_),
    .B1(_03854_),
    .B2(_06294_),
    .ZN(_06322_));
 OR2_X1 _23400_ (.A1(_06321_),
    .A2(_06322_),
    .ZN(_01272_));
 AOI21_X1 _23401_ (.A(_03927_),
    .B1(_03881_),
    .B2(_03478_),
    .ZN(_01273_));
 OAI22_X1 _23402_ (.A1(_03947_),
    .A2(_03873_),
    .B1(_03924_),
    .B2(_03918_),
    .ZN(_01274_));
 AOI21_X1 _23403_ (.A(net309),
    .B1(_05314_),
    .B2(_05338_),
    .ZN(_06323_));
 NAND2_X1 _23404_ (.A1(_10909_),
    .A2(_06261_),
    .ZN(_06324_));
 OAI21_X1 _23405_ (.A(_03439_),
    .B1(_06323_),
    .B2(_06324_),
    .ZN(_06325_));
 AOI22_X1 _23406_ (.A1(_06257_),
    .A2(_06258_),
    .B1(_06325_),
    .B2(_10350_),
    .ZN(_01275_));
 NAND2_X1 _23407_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .A2(_03613_),
    .ZN(_06326_));
 MUX2_X1 _23408_ (.A(_14068_),
    .B(_03660_),
    .S(_03780_),
    .Z(_06327_));
 OAI21_X1 _23409_ (.A(_06326_),
    .B1(_06327_),
    .B2(_03613_),
    .ZN(_01276_));
 NAND2_X1 _23410_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .A2(_03613_),
    .ZN(_06328_));
 MUX2_X1 _23411_ (.A(_05328_),
    .B(_11313_),
    .S(_03780_),
    .Z(_06329_));
 OAI21_X1 _23412_ (.A(_06328_),
    .B1(_06329_),
    .B2(_03613_),
    .ZN(_01277_));
 MUX2_X1 _23413_ (.A(\alu_adder_result_ex[11] ),
    .B(_11351_),
    .S(_03780_),
    .Z(_06330_));
 MUX2_X1 _23414_ (.A(_06330_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .S(_03613_),
    .Z(_01278_));
 MUX2_X1 _23415_ (.A(\alu_adder_result_ex[12] ),
    .B(_11993_),
    .S(_03780_),
    .Z(_06331_));
 CLKBUF_X3 _23416_ (.A(_03612_),
    .Z(_06332_));
 MUX2_X1 _23417_ (.A(_06331_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .S(_06332_),
    .Z(_01279_));
 MUX2_X1 _23418_ (.A(\alu_adder_result_ex[13] ),
    .B(_12044_),
    .S(_03780_),
    .Z(_06333_));
 MUX2_X1 _23419_ (.A(_06333_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .S(_06332_),
    .Z(_01280_));
 MUX2_X1 _23420_ (.A(net380),
    .B(_12144_),
    .S(_03780_),
    .Z(_06334_));
 MUX2_X1 _23421_ (.A(_06334_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .S(_06332_),
    .Z(_01281_));
 CLKBUF_X3 _23422_ (.A(_03779_),
    .Z(_06335_));
 MUX2_X1 _23423_ (.A(\alu_adder_result_ex[15] ),
    .B(_12221_),
    .S(_06335_),
    .Z(_06336_));
 MUX2_X1 _23424_ (.A(_06336_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .S(_06332_),
    .Z(_01282_));
 MUX2_X1 _23425_ (.A(\alu_adder_result_ex[16] ),
    .B(_12316_),
    .S(_06335_),
    .Z(_06337_));
 MUX2_X1 _23426_ (.A(_06337_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .S(_06332_),
    .Z(_01283_));
 MUX2_X1 _23427_ (.A(\alu_adder_result_ex[17] ),
    .B(net344),
    .S(_06335_),
    .Z(_06338_));
 MUX2_X1 _23428_ (.A(_06338_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .S(_06332_),
    .Z(_01284_));
 MUX2_X1 _23429_ (.A(net370),
    .B(net347),
    .S(_06335_),
    .Z(_06339_));
 MUX2_X1 _23430_ (.A(_06339_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .S(_06332_),
    .Z(_01285_));
 MUX2_X1 _23431_ (.A(net381),
    .B(net349),
    .S(_06335_),
    .Z(_06340_));
 MUX2_X1 _23432_ (.A(_06340_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .S(_06332_),
    .Z(_01286_));
 MUX2_X1 _23433_ (.A(\alu_adder_result_ex[1] ),
    .B(net348),
    .S(_06335_),
    .Z(_06341_));
 MUX2_X1 _23434_ (.A(_06341_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .S(_06332_),
    .Z(_01287_));
 MUX2_X1 _23435_ (.A(\alu_adder_result_ex[20] ),
    .B(_12651_),
    .S(_06335_),
    .Z(_06342_));
 MUX2_X1 _23436_ (.A(_06342_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .S(_06332_),
    .Z(_01288_));
 MUX2_X1 _23437_ (.A(net366),
    .B(_12725_),
    .S(_06335_),
    .Z(_06343_));
 CLKBUF_X3 _23438_ (.A(_03612_),
    .Z(_06344_));
 MUX2_X1 _23439_ (.A(_06343_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .S(_06344_),
    .Z(_01289_));
 MUX2_X1 _23440_ (.A(\alu_adder_result_ex[22] ),
    .B(_12823_),
    .S(_06335_),
    .Z(_06345_));
 MUX2_X1 _23441_ (.A(_06345_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .S(_06344_),
    .Z(_01290_));
 MUX2_X1 _23442_ (.A(net372),
    .B(net285),
    .S(_06335_),
    .Z(_06346_));
 MUX2_X1 _23443_ (.A(_06346_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .S(_06344_),
    .Z(_01291_));
 CLKBUF_X3 _23444_ (.A(_03779_),
    .Z(_06347_));
 MUX2_X1 _23445_ (.A(\alu_adder_result_ex[24] ),
    .B(_12985_),
    .S(_06347_),
    .Z(_06348_));
 MUX2_X1 _23446_ (.A(_06348_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .S(_06344_),
    .Z(_01292_));
 MUX2_X1 _23447_ (.A(net373),
    .B(net292),
    .S(_06347_),
    .Z(_06349_));
 MUX2_X1 _23448_ (.A(_06349_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .S(_06344_),
    .Z(_01293_));
 MUX2_X1 _23449_ (.A(net383),
    .B(_13155_),
    .S(_06347_),
    .Z(_06350_));
 MUX2_X1 _23450_ (.A(_06350_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .S(_06344_),
    .Z(_01294_));
 MUX2_X1 _23451_ (.A(net376),
    .B(_13224_),
    .S(_06347_),
    .Z(_06351_));
 MUX2_X1 _23452_ (.A(_06351_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .S(_06344_),
    .Z(_01295_));
 MUX2_X1 _23453_ (.A(\alu_adder_result_ex[28] ),
    .B(_13314_),
    .S(_06347_),
    .Z(_06352_));
 MUX2_X1 _23454_ (.A(_06352_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .S(_06344_),
    .Z(_01296_));
 MUX2_X1 _23455_ (.A(net14),
    .B(_03166_),
    .S(_06347_),
    .Z(_06353_));
 MUX2_X1 _23456_ (.A(_06353_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .S(_06344_),
    .Z(_01297_));
 MUX2_X1 _23457_ (.A(\alu_adder_result_ex[2] ),
    .B(_10973_),
    .S(_06347_),
    .Z(_06354_));
 MUX2_X1 _23458_ (.A(_06354_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .S(_06344_),
    .Z(_01298_));
 MUX2_X1 _23459_ (.A(\alu_adder_result_ex[30] ),
    .B(_03275_),
    .S(_06347_),
    .Z(_06355_));
 MUX2_X1 _23460_ (.A(_06355_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .S(_03612_),
    .Z(_01299_));
 NAND2_X1 _23461_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .A2(_03613_),
    .ZN(_06356_));
 OAI21_X1 _23462_ (.A(_03772_),
    .B1(net279),
    .B2(_03780_),
    .ZN(_06357_));
 OAI21_X1 _23463_ (.A(_06356_),
    .B1(_06357_),
    .B2(_03613_),
    .ZN(_01300_));
 NAND4_X2 _23464_ (.A1(_10310_),
    .A2(_10380_),
    .A3(_10873_),
    .A4(_10917_),
    .ZN(_06358_));
 NAND2_X1 _23465_ (.A1(_03790_),
    .A2(_06358_),
    .ZN(_06359_));
 NAND2_X1 _23466_ (.A1(_03650_),
    .A2(_06359_),
    .ZN(_06360_));
 NOR3_X1 _23467_ (.A1(_03779_),
    .A2(_03790_),
    .A3(_06358_),
    .ZN(_06361_));
 AOI21_X1 _23468_ (.A(_06361_),
    .B1(_03790_),
    .B2(_03779_),
    .ZN(_06362_));
 AOI21_X4 _23469_ (.A(_10912_),
    .B1(_10526_),
    .B2(_10874_),
    .ZN(_06363_));
 AOI21_X1 _23470_ (.A(_06362_),
    .B1(_06363_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .ZN(_06364_));
 INV_X1 _23471_ (.A(_03611_),
    .ZN(_06365_));
 NAND3_X4 _23472_ (.A1(_03407_),
    .A2(_06365_),
    .A3(_04033_),
    .ZN(_06366_));
 OAI22_X1 _23473_ (.A1(_06360_),
    .A2(_06364_),
    .B1(_06366_),
    .B2(_03647_),
    .ZN(_06367_));
 AND2_X1 _23474_ (.A1(_10310_),
    .A2(_06367_),
    .ZN(_06368_));
 NOR3_X1 _23475_ (.A1(_11408_),
    .A2(_11428_),
    .A3(_06368_),
    .ZN(_06369_));
 CLKBUF_X3 _23476_ (.A(_06369_),
    .Z(_06370_));
 CLKBUF_X3 _23477_ (.A(_06370_),
    .Z(_06371_));
 NAND2_X1 _23478_ (.A1(_05349_),
    .A2(_06371_),
    .ZN(_06372_));
 OR3_X1 _23479_ (.A1(_11406_),
    .A2(_11428_),
    .A3(_06368_),
    .ZN(_06373_));
 CLKBUF_X3 _23480_ (.A(_06373_),
    .Z(_06374_));
 NOR2_X2 _23481_ (.A1(_03450_),
    .A2(_06374_),
    .ZN(_06375_));
 NOR4_X4 _23482_ (.A1(_11432_),
    .A2(_10488_),
    .A3(_10508_),
    .A4(_10541_),
    .ZN(_06376_));
 AND2_X1 _23483_ (.A1(_06376_),
    .A2(_06363_),
    .ZN(_06377_));
 BUF_X4 _23484_ (.A(_06377_),
    .Z(_06378_));
 NOR2_X2 _23485_ (.A1(_06366_),
    .A2(_06378_),
    .ZN(_06379_));
 NAND2_X1 _23486_ (.A1(_06375_),
    .A2(_06379_),
    .ZN(_06380_));
 BUF_X4 _23487_ (.A(_06380_),
    .Z(_06381_));
 BUF_X4 _23488_ (.A(_06381_),
    .Z(_06382_));
 CLKBUF_X3 _23489_ (.A(_06370_),
    .Z(_06383_));
 OAI221_X1 _23490_ (.A(_06372_),
    .B1(_06382_),
    .B2(_04045_),
    .C1(_06383_),
    .C2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .ZN(_06384_));
 CLKBUF_X3 _23491_ (.A(_03404_),
    .Z(_06385_));
 CLKBUF_X3 _23492_ (.A(_06385_),
    .Z(_06386_));
 CLKBUF_X3 _23493_ (.A(_06378_),
    .Z(_06387_));
 XOR2_X2 _23494_ (.A(_03408_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .Z(_06388_));
 NAND2_X2 _23495_ (.A1(_03412_),
    .A2(_06388_),
    .ZN(_06389_));
 OAI21_X4 _23496_ (.A(_06389_),
    .B1(_06388_),
    .B2(net275),
    .ZN(_06390_));
 CLKBUF_X3 _23497_ (.A(_06390_),
    .Z(_06391_));
 BUF_X4 _23498_ (.A(_06391_),
    .Z(_06392_));
 MUX2_X1 _23499_ (.A(_14068_),
    .B(_00217_),
    .S(_06392_),
    .Z(_06393_));
 NOR2_X1 _23500_ (.A1(_06387_),
    .A2(_06393_),
    .ZN(_06394_));
 NAND2_X4 _23501_ (.A1(_06376_),
    .A2(_06363_),
    .ZN(_06395_));
 CLKBUF_X3 _23502_ (.A(_06395_),
    .Z(_06396_));
 CLKBUF_X3 _23503_ (.A(_06396_),
    .Z(_06397_));
 NAND2_X1 _23504_ (.A1(_03442_),
    .A2(_15540_),
    .ZN(_06398_));
 BUF_X4 _23505_ (.A(_06390_),
    .Z(_06399_));
 OR3_X2 _23506_ (.A1(_03444_),
    .A2(_03445_),
    .A3(_06399_),
    .ZN(_06400_));
 OR2_X1 _23507_ (.A1(_06398_),
    .A2(_06400_),
    .ZN(_06401_));
 AND2_X1 _23508_ (.A1(_00068_),
    .A2(_06401_),
    .ZN(_06402_));
 NOR2_X1 _23509_ (.A1(_06397_),
    .A2(_06402_),
    .ZN(_06403_));
 OAI21_X1 _23510_ (.A(_06386_),
    .B1(_06394_),
    .B2(_06403_),
    .ZN(_06404_));
 NAND2_X2 _23511_ (.A1(_06366_),
    .A2(_06375_),
    .ZN(_06405_));
 BUF_X4 _23512_ (.A(_06405_),
    .Z(_06406_));
 BUF_X4 _23513_ (.A(_06406_),
    .Z(_06407_));
 INV_X1 _23514_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .ZN(_06408_));
 CLKBUF_X3 _23515_ (.A(_15541_),
    .Z(_06409_));
 MUX2_X1 _23516_ (.A(_00118_),
    .B(_00116_),
    .S(_06409_),
    .Z(_06410_));
 MUX2_X1 _23517_ (.A(_00119_),
    .B(_00117_),
    .S(_06409_),
    .Z(_06411_));
 BUF_X4 _23518_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_06412_));
 MUX2_X1 _23519_ (.A(_06410_),
    .B(_06411_),
    .S(_06412_),
    .Z(_06413_));
 MUX2_X1 _23520_ (.A(_00126_),
    .B(_00124_),
    .S(_06409_),
    .Z(_06414_));
 MUX2_X1 _23521_ (.A(_00127_),
    .B(_00125_),
    .S(_06409_),
    .Z(_06415_));
 MUX2_X1 _23522_ (.A(_06414_),
    .B(_06415_),
    .S(_06412_),
    .Z(_06416_));
 NOR3_X2 _23523_ (.A1(_03445_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A3(_06412_),
    .ZN(_06417_));
 XNOR2_X2 _23524_ (.A(_00067_),
    .B(_06417_),
    .ZN(_06418_));
 MUX2_X1 _23525_ (.A(_06413_),
    .B(_06416_),
    .S(_06418_),
    .Z(_06419_));
 MUX2_X1 _23526_ (.A(_00122_),
    .B(_00120_),
    .S(_06409_),
    .Z(_06420_));
 BUF_X4 _23527_ (.A(_06409_),
    .Z(_06421_));
 MUX2_X1 _23528_ (.A(_00123_),
    .B(_00121_),
    .S(_06421_),
    .Z(_06422_));
 MUX2_X1 _23529_ (.A(_06420_),
    .B(_06422_),
    .S(_06412_),
    .Z(_06423_));
 MUX2_X1 _23530_ (.A(_00130_),
    .B(_00128_),
    .S(_06409_),
    .Z(_06424_));
 MUX2_X1 _23531_ (.A(_00131_),
    .B(_00129_),
    .S(_06421_),
    .Z(_06425_));
 MUX2_X1 _23532_ (.A(_06424_),
    .B(_06425_),
    .S(_06412_),
    .Z(_06426_));
 MUX2_X1 _23533_ (.A(_06423_),
    .B(_06426_),
    .S(_06418_),
    .Z(_06427_));
 XNOR2_X2 _23534_ (.A(_15542_),
    .B(_00066_),
    .ZN(_06428_));
 MUX2_X1 _23535_ (.A(_06419_),
    .B(_06427_),
    .S(_06428_),
    .Z(_06429_));
 MUX2_X1 _23536_ (.A(_00102_),
    .B(_00100_),
    .S(_06409_),
    .Z(_06430_));
 MUX2_X1 _23537_ (.A(_00103_),
    .B(_00101_),
    .S(_06421_),
    .Z(_06431_));
 MUX2_X1 _23538_ (.A(_06430_),
    .B(_06431_),
    .S(_06412_),
    .Z(_06432_));
 MUX2_X1 _23539_ (.A(_00110_),
    .B(_00108_),
    .S(_06421_),
    .Z(_06433_));
 MUX2_X1 _23540_ (.A(_00111_),
    .B(_00109_),
    .S(_06421_),
    .Z(_06434_));
 MUX2_X1 _23541_ (.A(_06433_),
    .B(_06434_),
    .S(_06412_),
    .Z(_06435_));
 MUX2_X1 _23542_ (.A(_06432_),
    .B(_06435_),
    .S(_06418_),
    .Z(_06436_));
 MUX2_X1 _23543_ (.A(_00106_),
    .B(_00104_),
    .S(_06421_),
    .Z(_06437_));
 MUX2_X1 _23544_ (.A(_00107_),
    .B(_00105_),
    .S(_06421_),
    .Z(_06438_));
 MUX2_X1 _23545_ (.A(_06437_),
    .B(_06438_),
    .S(_06412_),
    .Z(_06439_));
 MUX2_X1 _23546_ (.A(_00114_),
    .B(_00112_),
    .S(_06421_),
    .Z(_06440_));
 MUX2_X1 _23547_ (.A(_00115_),
    .B(_00113_),
    .S(_06421_),
    .Z(_06441_));
 MUX2_X1 _23548_ (.A(_06440_),
    .B(_06441_),
    .S(_06412_),
    .Z(_06442_));
 MUX2_X1 _23549_ (.A(_06439_),
    .B(_06442_),
    .S(_06418_),
    .Z(_06443_));
 MUX2_X1 _23550_ (.A(_06436_),
    .B(_06443_),
    .S(_06428_),
    .Z(_06444_));
 NAND2_X1 _23551_ (.A1(_15542_),
    .A2(_03446_),
    .ZN(_06445_));
 XNOR2_X2 _23552_ (.A(_03442_),
    .B(_06445_),
    .ZN(_06446_));
 MUX2_X1 _23553_ (.A(_06429_),
    .B(_06444_),
    .S(_06446_),
    .Z(_06447_));
 OAI222_X2 _23554_ (.A1(_03401_),
    .A2(_14068_),
    .B1(_06408_),
    .B2(_06365_),
    .C1(_06447_),
    .C2(_03432_),
    .ZN(_06448_));
 NOR2_X1 _23555_ (.A1(_06407_),
    .A2(_06448_),
    .ZN(_06449_));
 AOI21_X1 _23556_ (.A(_06384_),
    .B1(_06404_),
    .B2(_06449_),
    .ZN(_01301_));
 CLKBUF_X3 _23557_ (.A(_06374_),
    .Z(_06450_));
 NAND2_X1 _23558_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_06450_),
    .ZN(_06451_));
 NOR4_X4 _23559_ (.A1(_03403_),
    .A2(_03404_),
    .A3(_03650_),
    .A4(_03611_),
    .ZN(_06452_));
 BUF_X4 _23560_ (.A(_06452_),
    .Z(_06453_));
 NOR2_X1 _23561_ (.A1(_03450_),
    .A2(_06453_),
    .ZN(_06454_));
 OAI221_X1 _23562_ (.A(_06454_),
    .B1(_16090_),
    .B2(_03401_),
    .C1(_03432_),
    .C2(_06393_),
    .ZN(_06455_));
 CLKBUF_X3 _23563_ (.A(_06391_),
    .Z(_06456_));
 NOR2_X1 _23564_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_06456_),
    .ZN(_06457_));
 AOI21_X2 _23565_ (.A(_06457_),
    .B1(_06392_),
    .B2(_00185_),
    .ZN(_06458_));
 NOR2_X1 _23566_ (.A1(_06387_),
    .A2(_06458_),
    .ZN(_06459_));
 INV_X1 _23567_ (.A(_00069_),
    .ZN(_06460_));
 NOR3_X2 _23568_ (.A1(_03444_),
    .A2(_03445_),
    .A3(_06392_),
    .ZN(_06461_));
 AOI21_X2 _23569_ (.A(_06460_),
    .B1(_03443_),
    .B2(_06461_),
    .ZN(_06462_));
 AOI21_X1 _23570_ (.A(_06459_),
    .B1(_06462_),
    .B2(_06387_),
    .ZN(_06463_));
 AOI21_X1 _23571_ (.A(_06455_),
    .B1(_06463_),
    .B2(_06386_),
    .ZN(_06464_));
 NAND2_X1 _23572_ (.A1(_03440_),
    .A2(_06379_),
    .ZN(_06465_));
 OAI221_X1 _23573_ (.A(_06383_),
    .B1(_06465_),
    .B2(_03681_),
    .C1(_05389_),
    .C2(_10495_),
    .ZN(_06466_));
 OAI21_X1 _23574_ (.A(_06451_),
    .B1(_06464_),
    .B2(_06466_),
    .ZN(_01302_));
 NAND2_X1 _23575_ (.A1(_05431_),
    .A2(_06374_),
    .ZN(_06467_));
 OAI221_X1 _23576_ (.A(_06467_),
    .B1(_06450_),
    .B2(_05430_),
    .C1(net293),
    .C2(_06382_),
    .ZN(_06468_));
 CLKBUF_X3 _23577_ (.A(_06385_),
    .Z(_06469_));
 NAND2_X1 _23578_ (.A1(_03442_),
    .A2(_15544_),
    .ZN(_06470_));
 OAI21_X1 _23579_ (.A(_00070_),
    .B1(_06400_),
    .B2(_06470_),
    .ZN(_06471_));
 NOR2_X1 _23580_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_06456_),
    .ZN(_06472_));
 BUF_X4 _23581_ (.A(_06399_),
    .Z(_06473_));
 CLKBUF_X3 _23582_ (.A(_06473_),
    .Z(_06474_));
 AOI21_X1 _23583_ (.A(_06472_),
    .B1(_06474_),
    .B2(_00556_),
    .ZN(_06475_));
 MUX2_X1 _23584_ (.A(_06471_),
    .B(_06475_),
    .S(_06397_),
    .Z(_06476_));
 NAND2_X1 _23585_ (.A1(_06469_),
    .A2(_06476_),
    .ZN(_06477_));
 BUF_X4 _23586_ (.A(_03431_),
    .Z(_06478_));
 INV_X2 _23587_ (.A(_03401_),
    .ZN(_06479_));
 AOI221_X2 _23588_ (.A(_06407_),
    .B1(_06458_),
    .B2(_06478_),
    .C1(_06479_),
    .C2(\alu_adder_result_ex[2] ),
    .ZN(_06480_));
 AOI21_X1 _23589_ (.A(_06468_),
    .B1(_06477_),
    .B2(_06480_),
    .ZN(_01303_));
 NAND2_X1 _23590_ (.A1(_05469_),
    .A2(_06371_),
    .ZN(_06481_));
 BUF_X4 _23591_ (.A(_06370_),
    .Z(_06482_));
 OAI221_X1 _23592_ (.A(_06481_),
    .B1(_06382_),
    .B2(net319),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .C2(_06482_),
    .ZN(_06483_));
 NAND2_X2 _23593_ (.A1(_03442_),
    .A2(_15548_),
    .ZN(_06484_));
 OAI21_X1 _23594_ (.A(_00071_),
    .B1(_06400_),
    .B2(_06484_),
    .ZN(_06485_));
 NOR2_X1 _23595_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_06392_),
    .ZN(_06486_));
 AOI21_X1 _23596_ (.A(_06486_),
    .B1(_06474_),
    .B2(_00557_),
    .ZN(_06487_));
 MUX2_X1 _23597_ (.A(_06485_),
    .B(_06487_),
    .S(_06397_),
    .Z(_06488_));
 NAND2_X1 _23598_ (.A1(_06469_),
    .A2(_06488_),
    .ZN(_06489_));
 AOI221_X1 _23599_ (.A(_06407_),
    .B1(_06475_),
    .B2(_06478_),
    .C1(_06479_),
    .C2(\alu_adder_result_ex[3] ),
    .ZN(_06490_));
 AOI21_X1 _23600_ (.A(_06483_),
    .B1(_06489_),
    .B2(_06490_),
    .ZN(_01304_));
 NAND2_X1 _23601_ (.A1(_05523_),
    .A2(_06371_),
    .ZN(_06491_));
 OAI221_X2 _23602_ (.A(_06491_),
    .B1(_06382_),
    .B2(_11591_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .C2(_06482_),
    .ZN(_06492_));
 AOI221_X2 _23603_ (.A(_06407_),
    .B1(_06487_),
    .B2(_03614_),
    .C1(_06479_),
    .C2(\alu_adder_result_ex[4] ),
    .ZN(_06493_));
 OR3_X1 _23604_ (.A1(_03444_),
    .A2(_00066_),
    .A3(_06390_),
    .ZN(_06494_));
 BUF_X2 _23605_ (.A(_06494_),
    .Z(_06495_));
 OAI21_X1 _23606_ (.A(_00072_),
    .B1(_06398_),
    .B2(_06495_),
    .ZN(_06496_));
 NOR2_X1 _23607_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_06392_),
    .ZN(_06497_));
 AOI21_X1 _23608_ (.A(_06497_),
    .B1(_06474_),
    .B2(_00558_),
    .ZN(_06498_));
 MUX2_X1 _23609_ (.A(_06496_),
    .B(_06498_),
    .S(_06396_),
    .Z(_06499_));
 NAND2_X1 _23610_ (.A1(_06386_),
    .A2(_06499_),
    .ZN(_06500_));
 AOI21_X1 _23611_ (.A(_06492_),
    .B1(_06493_),
    .B2(_06500_),
    .ZN(_01305_));
 CLKBUF_X3 _23612_ (.A(_06369_),
    .Z(_06501_));
 NAND2_X1 _23613_ (.A1(_05556_),
    .A2(_06501_),
    .ZN(_06502_));
 OAI221_X2 _23614_ (.A(_06502_),
    .B1(_06382_),
    .B2(_11629_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .C2(_06482_),
    .ZN(_06503_));
 AOI221_X1 _23615_ (.A(_06407_),
    .B1(_06498_),
    .B2(_03614_),
    .C1(_06479_),
    .C2(\alu_adder_result_ex[5] ),
    .ZN(_06504_));
 NAND2_X1 _23616_ (.A1(_03442_),
    .A2(_15546_),
    .ZN(_06505_));
 OAI21_X1 _23617_ (.A(_00073_),
    .B1(_06505_),
    .B2(_06495_),
    .ZN(_06506_));
 NOR2_X1 _23618_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_06456_),
    .ZN(_06507_));
 AOI21_X1 _23619_ (.A(_06507_),
    .B1(_06474_),
    .B2(_00559_),
    .ZN(_06508_));
 MUX2_X1 _23620_ (.A(_06506_),
    .B(_06508_),
    .S(_06396_),
    .Z(_06509_));
 NAND2_X1 _23621_ (.A1(_06386_),
    .A2(_06509_),
    .ZN(_06510_));
 AOI21_X1 _23622_ (.A(_06503_),
    .B1(_06504_),
    .B2(_06510_),
    .ZN(_01306_));
 MUX2_X1 _23623_ (.A(\alu_adder_result_ex[3] ),
    .B(_11019_),
    .S(_06347_),
    .Z(_06511_));
 MUX2_X1 _23624_ (.A(_06511_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .S(_03612_),
    .Z(_01307_));
 NAND2_X1 _23625_ (.A1(_05591_),
    .A2(_06501_),
    .ZN(_06512_));
 OAI221_X2 _23626_ (.A(_06512_),
    .B1(_06382_),
    .B2(_11672_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .C2(_06482_),
    .ZN(_06513_));
 AOI221_X1 _23627_ (.A(_06407_),
    .B1(_06508_),
    .B2(_03614_),
    .C1(_06479_),
    .C2(\alu_adder_result_ex[6] ),
    .ZN(_06514_));
 OAI21_X1 _23628_ (.A(_00074_),
    .B1(_06470_),
    .B2(_06495_),
    .ZN(_06515_));
 NOR2_X1 _23629_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_06456_),
    .ZN(_06516_));
 AOI21_X1 _23630_ (.A(_06516_),
    .B1(_06474_),
    .B2(_00560_),
    .ZN(_06517_));
 MUX2_X1 _23631_ (.A(_06515_),
    .B(_06517_),
    .S(_06396_),
    .Z(_06518_));
 NAND2_X1 _23632_ (.A1(_06386_),
    .A2(_06518_),
    .ZN(_06519_));
 AOI21_X1 _23633_ (.A(_06513_),
    .B1(_06514_),
    .B2(_06519_),
    .ZN(_01308_));
 NAND2_X1 _23634_ (.A1(_05648_),
    .A2(_06501_),
    .ZN(_06520_));
 OAI221_X2 _23635_ (.A(_06520_),
    .B1(_06382_),
    .B2(_03723_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .C2(_06482_),
    .ZN(_06521_));
 AOI221_X2 _23636_ (.A(_06407_),
    .B1(_06517_),
    .B2(_03614_),
    .C1(_03652_),
    .C2(\alu_adder_result_ex[7] ),
    .ZN(_06522_));
 OAI21_X1 _23637_ (.A(_00075_),
    .B1(_06484_),
    .B2(_06495_),
    .ZN(_06523_));
 NOR2_X1 _23638_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_06456_),
    .ZN(_06524_));
 AOI21_X1 _23639_ (.A(_06524_),
    .B1(_06474_),
    .B2(_00561_),
    .ZN(_06525_));
 MUX2_X1 _23640_ (.A(_06523_),
    .B(_06525_),
    .S(_06396_),
    .Z(_06526_));
 NAND2_X1 _23641_ (.A1(_06386_),
    .A2(_06526_),
    .ZN(_06527_));
 AOI21_X1 _23642_ (.A(_06521_),
    .B1(_06522_),
    .B2(_06527_),
    .ZN(_01309_));
 NAND2_X1 _23643_ (.A1(_05664_),
    .A2(_06501_),
    .ZN(_06528_));
 OAI221_X1 _23644_ (.A(_06528_),
    .B1(_06381_),
    .B2(_03732_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .C2(_06482_),
    .ZN(_06529_));
 NOR2_X1 _23645_ (.A1(_03445_),
    .A2(_00067_),
    .ZN(_06530_));
 OAI211_X4 _23646_ (.A(_06389_),
    .B(_06530_),
    .C1(net276),
    .C2(_06388_),
    .ZN(_06531_));
 OAI21_X1 _23647_ (.A(_00076_),
    .B1(_06398_),
    .B2(_06531_),
    .ZN(_06532_));
 NOR2_X1 _23648_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_06456_),
    .ZN(_06533_));
 AOI21_X1 _23649_ (.A(_06533_),
    .B1(_06474_),
    .B2(_00562_),
    .ZN(_06534_));
 MUX2_X1 _23650_ (.A(_06532_),
    .B(_06534_),
    .S(_06397_),
    .Z(_06535_));
 NAND2_X1 _23651_ (.A1(_06469_),
    .A2(_06535_),
    .ZN(_06536_));
 AOI221_X2 _23652_ (.A(_06407_),
    .B1(_06525_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(\alu_adder_result_ex[8] ),
    .ZN(_06537_));
 AOI21_X1 _23653_ (.A(_06529_),
    .B1(_06536_),
    .B2(_06537_),
    .ZN(_01310_));
 NAND2_X1 _23654_ (.A1(_05700_),
    .A2(_06501_),
    .ZN(_06538_));
 OAI221_X1 _23655_ (.A(_06538_),
    .B1(_06381_),
    .B2(_11824_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .C2(_06482_),
    .ZN(_06539_));
 NOR2_X1 _23656_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_06473_),
    .ZN(_06540_));
 AOI21_X2 _23657_ (.A(_06540_),
    .B1(_06392_),
    .B2(_00563_),
    .ZN(_06541_));
 NOR2_X1 _23658_ (.A1(_06387_),
    .A2(_06541_),
    .ZN(_06542_));
 INV_X1 _23659_ (.A(_00077_),
    .ZN(_06543_));
 NOR3_X2 _23660_ (.A1(_03445_),
    .A2(_00067_),
    .A3(_06392_),
    .ZN(_06544_));
 AOI21_X2 _23661_ (.A(_06543_),
    .B1(_03443_),
    .B2(_06544_),
    .ZN(_06545_));
 AOI21_X1 _23662_ (.A(_06542_),
    .B1(_06545_),
    .B2(_06387_),
    .ZN(_06546_));
 NAND2_X1 _23663_ (.A1(_06469_),
    .A2(_06546_),
    .ZN(_06547_));
 AOI221_X2 _23664_ (.A(_06407_),
    .B1(_06534_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(\alu_adder_result_ex[9] ),
    .ZN(_06548_));
 AOI21_X1 _23665_ (.A(_06539_),
    .B1(_06547_),
    .B2(_06548_),
    .ZN(_01311_));
 NAND2_X1 _23666_ (.A1(_05724_),
    .A2(_06374_),
    .ZN(_06549_));
 OAI221_X1 _23667_ (.A(_06549_),
    .B1(_06450_),
    .B2(_05723_),
    .C1(_11898_),
    .C2(_06382_),
    .ZN(_06550_));
 OAI21_X1 _23668_ (.A(_00078_),
    .B1(_06470_),
    .B2(_06531_),
    .ZN(_06551_));
 NOR2_X1 _23669_ (.A1(net386),
    .A2(_06390_),
    .ZN(_06552_));
 AOI21_X1 _23670_ (.A(_06552_),
    .B1(_06399_),
    .B2(_00564_),
    .ZN(_06553_));
 MUX2_X1 _23671_ (.A(_06551_),
    .B(_06553_),
    .S(_06397_),
    .Z(_06554_));
 NAND2_X1 _23672_ (.A1(_06469_),
    .A2(_06554_),
    .ZN(_06555_));
 AOI221_X2 _23673_ (.A(_06406_),
    .B1(_06541_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(net386),
    .ZN(_06556_));
 AOI21_X1 _23674_ (.A(_06550_),
    .B1(_06555_),
    .B2(_06556_),
    .ZN(_01312_));
 NOR2_X1 _23675_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .A2(_06370_),
    .ZN(_06557_));
 AOI221_X1 _23676_ (.A(_06452_),
    .B1(_06553_),
    .B2(_03403_),
    .C1(_03650_),
    .C2(\alu_adder_result_ex[11] ),
    .ZN(_06558_));
 OAI211_X2 _23677_ (.A(_00079_),
    .B(_06378_),
    .C1(_06484_),
    .C2(_06531_),
    .ZN(_06559_));
 NOR2_X1 _23678_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_06391_),
    .ZN(_06560_));
 AOI21_X2 _23679_ (.A(_06560_),
    .B1(_06473_),
    .B2(_00565_),
    .ZN(_06561_));
 OAI21_X1 _23680_ (.A(_06559_),
    .B1(_06561_),
    .B2(_06378_),
    .ZN(_06562_));
 OAI21_X1 _23681_ (.A(_06558_),
    .B1(_06562_),
    .B2(_03452_),
    .ZN(_06563_));
 NAND2_X2 _23682_ (.A1(_06453_),
    .A2(_06395_),
    .ZN(_06564_));
 OAI21_X1 _23683_ (.A(_06563_),
    .B1(_06564_),
    .B2(net365),
    .ZN(_06565_));
 AOI221_X1 _23684_ (.A(_06557_),
    .B1(_06565_),
    .B2(_06375_),
    .C1(_05771_),
    .C2(_06371_),
    .ZN(_01313_));
 OAI21_X1 _23685_ (.A(_05816_),
    .B1(_06465_),
    .B2(_10868_),
    .ZN(_06566_));
 NOR2_X1 _23686_ (.A1(_06374_),
    .A2(_06566_),
    .ZN(_06567_));
 AOI21_X1 _23687_ (.A(_06567_),
    .B1(_06450_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .ZN(_06568_));
 OR3_X1 _23688_ (.A1(_00066_),
    .A2(_00067_),
    .A3(_06390_),
    .ZN(_06569_));
 BUF_X2 _23689_ (.A(_06569_),
    .Z(_06570_));
 OAI21_X1 _23690_ (.A(_00080_),
    .B1(_06398_),
    .B2(_06570_),
    .ZN(_06571_));
 NOR2_X1 _23691_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_06456_),
    .ZN(_06572_));
 AOI21_X1 _23692_ (.A(_06572_),
    .B1(_06474_),
    .B2(_00566_),
    .ZN(_06573_));
 MUX2_X1 _23693_ (.A(_06571_),
    .B(_06573_),
    .S(_06397_),
    .Z(_06574_));
 NAND2_X1 _23694_ (.A1(_06469_),
    .A2(_06574_),
    .ZN(_06575_));
 AOI221_X2 _23695_ (.A(_06406_),
    .B1(_06561_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(\alu_adder_result_ex[12] ),
    .ZN(_06576_));
 AOI21_X1 _23696_ (.A(_06568_),
    .B1(_06575_),
    .B2(_06576_),
    .ZN(_01314_));
 NAND2_X1 _23697_ (.A1(_04023_),
    .A2(_04626_),
    .ZN(_06577_));
 OAI21_X1 _23698_ (.A(_06577_),
    .B1(_05104_),
    .B2(_04626_),
    .ZN(_06578_));
 NAND3_X1 _23699_ (.A1(_12103_),
    .A2(_06501_),
    .A3(_06578_),
    .ZN(_06579_));
 OAI221_X1 _23700_ (.A(_06579_),
    .B1(_06381_),
    .B2(_12075_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .C2(_06371_),
    .ZN(_06580_));
 OAI21_X1 _23701_ (.A(_00081_),
    .B1(_06505_),
    .B2(_06570_),
    .ZN(_06581_));
 NOR2_X1 _23702_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_06456_),
    .ZN(_06582_));
 AOI21_X1 _23703_ (.A(_06582_),
    .B1(_06474_),
    .B2(_04023_),
    .ZN(_06583_));
 MUX2_X1 _23704_ (.A(_06581_),
    .B(_06583_),
    .S(_06397_),
    .Z(_06584_));
 NAND2_X1 _23705_ (.A1(_06469_),
    .A2(_06584_),
    .ZN(_06585_));
 AOI221_X2 _23706_ (.A(_06406_),
    .B1(_06573_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(\alu_adder_result_ex[13] ),
    .ZN(_06586_));
 AOI21_X1 _23707_ (.A(_06580_),
    .B1(_06585_),
    .B2(_06586_),
    .ZN(_01315_));
 NAND2_X1 _23708_ (.A1(_04026_),
    .A2(_04626_),
    .ZN(_06587_));
 OAI21_X1 _23709_ (.A(_06587_),
    .B1(_05158_),
    .B2(_04626_),
    .ZN(_06588_));
 NAND3_X1 _23710_ (.A1(_12103_),
    .A2(_06501_),
    .A3(_06588_),
    .ZN(_06589_));
 OAI221_X1 _23711_ (.A(_06589_),
    .B1(_06381_),
    .B2(_12177_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .C2(_06371_),
    .ZN(_06590_));
 OAI21_X1 _23712_ (.A(_00082_),
    .B1(_06470_),
    .B2(_06570_),
    .ZN(_06591_));
 NOR2_X1 _23713_ (.A1(net380),
    .A2(_06391_),
    .ZN(_06592_));
 AOI21_X1 _23714_ (.A(_06592_),
    .B1(_06473_),
    .B2(_04026_),
    .ZN(_06593_));
 MUX2_X1 _23715_ (.A(_06591_),
    .B(_06593_),
    .S(_06397_),
    .Z(_06594_));
 NAND2_X1 _23716_ (.A1(_06469_),
    .A2(_06594_),
    .ZN(_06595_));
 AOI221_X2 _23717_ (.A(_06406_),
    .B1(_06583_),
    .B2(_06478_),
    .C1(_03652_),
    .C2(net380),
    .ZN(_06596_));
 AOI21_X1 _23718_ (.A(_06590_),
    .B1(_06595_),
    .B2(_06596_),
    .ZN(_01316_));
 OAI22_X1 _23719_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .A2(_06370_),
    .B1(_06381_),
    .B2(_12254_),
    .ZN(_06597_));
 NOR2_X2 _23720_ (.A1(_10495_),
    .A2(_06374_),
    .ZN(_06598_));
 MUX2_X1 _23721_ (.A(_00659_),
    .B(_05219_),
    .S(_04791_),
    .Z(_06599_));
 AOI221_X2 _23722_ (.A(_06406_),
    .B1(_06593_),
    .B2(_03431_),
    .C1(_03651_),
    .C2(\alu_adder_result_ex[15] ),
    .ZN(_06600_));
 OAI21_X1 _23723_ (.A(_00083_),
    .B1(_06484_),
    .B2(_06570_),
    .ZN(_06601_));
 NOR2_X1 _23724_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_06473_),
    .ZN(_06602_));
 AOI21_X1 _23725_ (.A(_06602_),
    .B1(_06392_),
    .B2(_00659_),
    .ZN(_06603_));
 MUX2_X1 _23726_ (.A(_06601_),
    .B(_06603_),
    .S(_06395_),
    .Z(_06604_));
 NAND2_X1 _23727_ (.A1(_06385_),
    .A2(_06604_),
    .ZN(_06605_));
 AOI221_X1 _23728_ (.A(_06597_),
    .B1(_06598_),
    .B2(_06599_),
    .C1(_06600_),
    .C2(_06605_),
    .ZN(_01317_));
 MUX2_X1 _23729_ (.A(\alu_adder_result_ex[4] ),
    .B(_03519_),
    .S(_06347_),
    .Z(_06606_));
 MUX2_X1 _23730_ (.A(_06606_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .S(_03612_),
    .Z(_01318_));
 OR2_X1 _23731_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A2(_06370_),
    .ZN(_06607_));
 OAI221_X1 _23732_ (.A(_06607_),
    .B1(_06374_),
    .B2(_05991_),
    .C1(_12350_),
    .C2(_06382_),
    .ZN(_06608_));
 NOR2_X1 _23733_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_06473_),
    .ZN(_06609_));
 AOI21_X1 _23734_ (.A(_06609_),
    .B1(_06392_),
    .B2(_03670_),
    .ZN(_06610_));
 NOR2_X1 _23735_ (.A1(_06387_),
    .A2(_06610_),
    .ZN(_06611_));
 INV_X1 _23736_ (.A(_00084_),
    .ZN(_06612_));
 CLKBUF_X2 _23737_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .Z(_06613_));
 AND2_X1 _23738_ (.A1(_06613_),
    .A2(_15540_),
    .ZN(_06614_));
 AOI21_X2 _23739_ (.A(_06612_),
    .B1(_06461_),
    .B2(_06614_),
    .ZN(_06615_));
 AOI21_X1 _23740_ (.A(_06611_),
    .B1(_06615_),
    .B2(_06387_),
    .ZN(_06616_));
 NAND2_X1 _23741_ (.A1(_06469_),
    .A2(_06616_),
    .ZN(_06617_));
 AOI221_X2 _23742_ (.A(_06406_),
    .B1(_06603_),
    .B2(_06478_),
    .C1(_03651_),
    .C2(\alu_adder_result_ex[16] ),
    .ZN(_06618_));
 AOI21_X1 _23743_ (.A(_06608_),
    .B1(_06617_),
    .B2(_06618_),
    .ZN(_01319_));
 OR2_X1 _23744_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A2(_06370_),
    .ZN(_06619_));
 OAI221_X2 _23745_ (.A(_06619_),
    .B1(_06374_),
    .B2(_06027_),
    .C1(_12425_),
    .C2(_06382_),
    .ZN(_06620_));
 NAND2_X1 _23746_ (.A1(_06613_),
    .A2(_15546_),
    .ZN(_06621_));
 OAI21_X1 _23747_ (.A(_00085_),
    .B1(_06400_),
    .B2(_06621_),
    .ZN(_06622_));
 NOR2_X1 _23748_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_06456_),
    .ZN(_06623_));
 AOI21_X1 _23749_ (.A(_06623_),
    .B1(_06474_),
    .B2(_03800_),
    .ZN(_06624_));
 MUX2_X1 _23750_ (.A(_06622_),
    .B(_06624_),
    .S(_06397_),
    .Z(_06625_));
 NAND2_X1 _23751_ (.A1(_06469_),
    .A2(_06625_),
    .ZN(_06626_));
 AOI221_X1 _23752_ (.A(_06406_),
    .B1(_06610_),
    .B2(_06478_),
    .C1(_03651_),
    .C2(\alu_adder_result_ex[17] ),
    .ZN(_06627_));
 AOI21_X1 _23753_ (.A(_06620_),
    .B1(_06626_),
    .B2(_06627_),
    .ZN(_01320_));
 NAND2_X1 _23754_ (.A1(_06082_),
    .A2(_06501_),
    .ZN(_06628_));
 OAI221_X2 _23755_ (.A(_06628_),
    .B1(_06381_),
    .B2(_12514_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .C2(_06371_),
    .ZN(_06629_));
 NAND2_X1 _23756_ (.A1(_06613_),
    .A2(_15544_),
    .ZN(_06630_));
 OAI21_X1 _23757_ (.A(_00086_),
    .B1(_06400_),
    .B2(_06630_),
    .ZN(_06631_));
 NOR2_X1 _23758_ (.A1(net369),
    .A2(_06456_),
    .ZN(_06632_));
 AOI21_X1 _23759_ (.A(_06632_),
    .B1(_06392_),
    .B2(_03804_),
    .ZN(_06633_));
 MUX2_X1 _23760_ (.A(_06631_),
    .B(_06633_),
    .S(_06397_),
    .Z(_06634_));
 NAND2_X1 _23761_ (.A1(_06386_),
    .A2(_06634_),
    .ZN(_06635_));
 AOI221_X2 _23762_ (.A(_06406_),
    .B1(_06624_),
    .B2(_03431_),
    .C1(_03651_),
    .C2(net369),
    .ZN(_06636_));
 AOI21_X1 _23763_ (.A(_06629_),
    .B1(_06635_),
    .B2(_06636_),
    .ZN(_01321_));
 NAND2_X1 _23764_ (.A1(_06111_),
    .A2(_06501_),
    .ZN(_06637_));
 OAI221_X1 _23765_ (.A(_06637_),
    .B1(_06381_),
    .B2(_12589_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .C2(_06371_),
    .ZN(_06638_));
 NAND2_X1 _23766_ (.A1(_06613_),
    .A2(_15548_),
    .ZN(_06639_));
 OAI21_X1 _23767_ (.A(_00087_),
    .B1(_06400_),
    .B2(_06639_),
    .ZN(_06640_));
 MUX2_X1 _23768_ (.A(net381),
    .B(_03806_),
    .S(_06399_),
    .Z(_06641_));
 MUX2_X1 _23769_ (.A(_06640_),
    .B(_06641_),
    .S(_06396_),
    .Z(_06642_));
 NAND2_X1 _23770_ (.A1(_06386_),
    .A2(_06642_),
    .ZN(_06643_));
 AOI221_X2 _23771_ (.A(_06406_),
    .B1(_06633_),
    .B2(_03431_),
    .C1(_03651_),
    .C2(net381),
    .ZN(_06644_));
 AOI21_X1 _23772_ (.A(_06638_),
    .B1(_06643_),
    .B2(_06644_),
    .ZN(_01322_));
 OAI22_X2 _23773_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_06370_),
    .B1(_06381_),
    .B2(net358),
    .ZN(_06645_));
 AOI221_X2 _23774_ (.A(_06405_),
    .B1(_06641_),
    .B2(_03403_),
    .C1(_03651_),
    .C2(\alu_adder_result_ex[20] ),
    .ZN(_06646_));
 NAND2_X1 _23775_ (.A1(_06613_),
    .A2(_15540_),
    .ZN(_06647_));
 OAI21_X1 _23776_ (.A(_00088_),
    .B1(_06495_),
    .B2(_06647_),
    .ZN(_06648_));
 NOR2_X1 _23777_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_06391_),
    .ZN(_06649_));
 AOI21_X1 _23778_ (.A(_06649_),
    .B1(_06473_),
    .B2(_03808_),
    .ZN(_06650_));
 MUX2_X1 _23779_ (.A(_06648_),
    .B(_06650_),
    .S(_06395_),
    .Z(_06651_));
 NAND2_X1 _23780_ (.A1(_06385_),
    .A2(_06651_),
    .ZN(_06652_));
 NOR2_X1 _23781_ (.A1(_10495_),
    .A2(_06154_),
    .ZN(_06653_));
 AOI221_X2 _23782_ (.A(_06645_),
    .B1(_06646_),
    .B2(_06652_),
    .C1(_06482_),
    .C2(_06653_),
    .ZN(_01323_));
 AND2_X1 _23783_ (.A1(_06182_),
    .A2(_06183_),
    .ZN(_06654_));
 NAND2_X1 _23784_ (.A1(_06654_),
    .A2(_06501_),
    .ZN(_06655_));
 OAI221_X1 _23785_ (.A(_06655_),
    .B1(_06381_),
    .B2(net363),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .C2(_06371_),
    .ZN(_06656_));
 AOI221_X2 _23786_ (.A(_06407_),
    .B1(_06650_),
    .B2(_03614_),
    .C1(_03652_),
    .C2(net366),
    .ZN(_06657_));
 OAI21_X1 _23787_ (.A(_00089_),
    .B1(_06495_),
    .B2(_06621_),
    .ZN(_06658_));
 MUX2_X1 _23788_ (.A(net366),
    .B(_03810_),
    .S(_06399_),
    .Z(_06659_));
 MUX2_X1 _23789_ (.A(_06658_),
    .B(_06659_),
    .S(_06396_),
    .Z(_06660_));
 NAND2_X1 _23790_ (.A1(_06386_),
    .A2(_06660_),
    .ZN(_06661_));
 AOI21_X1 _23791_ (.A(_06656_),
    .B1(_06657_),
    .B2(_06661_),
    .ZN(_01324_));
 NAND2_X1 _23792_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_06450_),
    .ZN(_06662_));
 AOI221_X2 _23793_ (.A(_06453_),
    .B1(_06659_),
    .B2(_03403_),
    .C1(_03650_),
    .C2(\alu_adder_result_ex[22] ),
    .ZN(_06663_));
 AOI21_X1 _23794_ (.A(_06663_),
    .B1(_06379_),
    .B2(_12859_),
    .ZN(_06664_));
 OAI21_X1 _23795_ (.A(_00090_),
    .B1(_06495_),
    .B2(_06630_),
    .ZN(_06665_));
 NOR2_X1 _23796_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_06399_),
    .ZN(_06666_));
 AOI21_X1 _23797_ (.A(_06666_),
    .B1(_06391_),
    .B2(_03813_),
    .ZN(_06667_));
 MUX2_X1 _23798_ (.A(_06665_),
    .B(_06667_),
    .S(_06396_),
    .Z(_06668_));
 AOI21_X1 _23799_ (.A(_06664_),
    .B1(_06668_),
    .B2(_06385_),
    .ZN(_06669_));
 NAND2_X1 _23800_ (.A1(_03440_),
    .A2(_06371_),
    .ZN(_06670_));
 INV_X1 _23801_ (.A(_06598_),
    .ZN(_06671_));
 OAI221_X1 _23802_ (.A(_06662_),
    .B1(_06669_),
    .B2(_06670_),
    .C1(_06671_),
    .C2(_04503_),
    .ZN(_01325_));
 OAI22_X1 _23803_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_06370_),
    .B1(_06380_),
    .B2(_03724_),
    .ZN(_06672_));
 AOI221_X2 _23804_ (.A(_06405_),
    .B1(_06667_),
    .B2(_03403_),
    .C1(_03651_),
    .C2(net372),
    .ZN(_06673_));
 OAI21_X1 _23805_ (.A(_00091_),
    .B1(_06495_),
    .B2(_06639_),
    .ZN(_06674_));
 NOR2_X1 _23806_ (.A1(net372),
    .A2(_06391_),
    .ZN(_06675_));
 AOI21_X2 _23807_ (.A(_06675_),
    .B1(_06473_),
    .B2(_03815_),
    .ZN(_06676_));
 MUX2_X1 _23808_ (.A(_06674_),
    .B(_06676_),
    .S(_06395_),
    .Z(_06677_));
 NAND2_X1 _23809_ (.A1(_06385_),
    .A2(_06677_),
    .ZN(_06678_));
 INV_X1 _23810_ (.A(_04659_),
    .ZN(_06679_));
 AOI221_X1 _23811_ (.A(_06672_),
    .B1(_06673_),
    .B2(_06678_),
    .C1(_06482_),
    .C2(_06679_),
    .ZN(_01326_));
 NAND2_X1 _23812_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(_06450_),
    .ZN(_06680_));
 AOI21_X1 _23813_ (.A(_06453_),
    .B1(\alu_adder_result_ex[24] ),
    .B2(_03650_),
    .ZN(_06681_));
 INV_X1 _23814_ (.A(_06681_),
    .ZN(_06682_));
 OAI21_X1 _23815_ (.A(_00092_),
    .B1(_06531_),
    .B2(_06647_),
    .ZN(_06683_));
 NOR2_X1 _23816_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_06399_),
    .ZN(_06684_));
 AOI21_X1 _23817_ (.A(_06684_),
    .B1(_06391_),
    .B2(_03817_),
    .ZN(_06685_));
 MUX2_X1 _23818_ (.A(_06683_),
    .B(_06685_),
    .S(_06395_),
    .Z(_06686_));
 AOI221_X2 _23819_ (.A(_06682_),
    .B1(_06686_),
    .B2(_03404_),
    .C1(_06676_),
    .C2(_03614_),
    .ZN(_06687_));
 AOI21_X1 _23820_ (.A(_03450_),
    .B1(_06379_),
    .B2(_13023_),
    .ZN(_06688_));
 NAND2_X1 _23821_ (.A1(_06482_),
    .A2(_06688_),
    .ZN(_06689_));
 OAI221_X1 _23822_ (.A(_06680_),
    .B1(_06687_),
    .B2(_06689_),
    .C1(_06671_),
    .C2(_04890_),
    .ZN(_01327_));
 AOI21_X1 _23823_ (.A(_06453_),
    .B1(net373),
    .B2(_03650_),
    .ZN(_06690_));
 INV_X1 _23824_ (.A(_06690_),
    .ZN(_06691_));
 OAI21_X1 _23825_ (.A(_00093_),
    .B1(_06531_),
    .B2(_06621_),
    .ZN(_06692_));
 NOR2_X1 _23826_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_06399_),
    .ZN(_06693_));
 AOI21_X1 _23827_ (.A(_06693_),
    .B1(_06391_),
    .B2(_03819_),
    .ZN(_06694_));
 MUX2_X1 _23828_ (.A(_06692_),
    .B(_06694_),
    .S(_06395_),
    .Z(_06695_));
 AOI221_X2 _23829_ (.A(_06691_),
    .B1(_06695_),
    .B2(_03404_),
    .C1(_06685_),
    .C2(_03431_),
    .ZN(_06696_));
 NOR2_X1 _23830_ (.A1(_13097_),
    .A2(_06564_),
    .ZN(_06697_));
 OAI21_X1 _23831_ (.A(_06375_),
    .B1(_06696_),
    .B2(_06697_),
    .ZN(_06698_));
 MUX2_X1 _23832_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B(_04949_),
    .S(_06370_),
    .Z(_06699_));
 AND2_X1 _23833_ (.A1(_06698_),
    .A2(_06699_),
    .ZN(_01328_));
 MUX2_X1 _23834_ (.A(\alu_adder_result_ex[5] ),
    .B(_03696_),
    .S(_03779_),
    .Z(_06700_));
 MUX2_X1 _23835_ (.A(_06700_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .S(_03612_),
    .Z(_01329_));
 AOI221_X1 _23836_ (.A(_06453_),
    .B1(_06694_),
    .B2(_03431_),
    .C1(_03651_),
    .C2(net382),
    .ZN(_06701_));
 OAI21_X1 _23837_ (.A(_00094_),
    .B1(_06531_),
    .B2(_06630_),
    .ZN(_06702_));
 MUX2_X1 _23838_ (.A(net382),
    .B(_03821_),
    .S(_06390_),
    .Z(_06703_));
 MUX2_X1 _23839_ (.A(_06702_),
    .B(_06703_),
    .S(_06395_),
    .Z(_06704_));
 NAND2_X1 _23840_ (.A1(_06385_),
    .A2(_06704_),
    .ZN(_06705_));
 NAND2_X1 _23841_ (.A1(_06701_),
    .A2(_06705_),
    .ZN(_06706_));
 OR2_X1 _23842_ (.A1(net352),
    .A2(_06564_),
    .ZN(_06707_));
 NAND4_X1 _23843_ (.A1(_03440_),
    .A2(_06383_),
    .A3(_06706_),
    .A4(_06707_),
    .ZN(_06708_));
 INV_X1 _23844_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .ZN(_06709_));
 OAI221_X1 _23845_ (.A(_06708_),
    .B1(_06671_),
    .B2(_05002_),
    .C1(_06709_),
    .C2(_06383_),
    .ZN(_01330_));
 AOI221_X2 _23846_ (.A(_06452_),
    .B1(_06703_),
    .B2(_03403_),
    .C1(_03650_),
    .C2(net377),
    .ZN(_06710_));
 OR2_X1 _23847_ (.A1(_06531_),
    .A2(_06639_),
    .ZN(_06711_));
 NAND3_X1 _23848_ (.A1(_00095_),
    .A2(_06378_),
    .A3(_06711_),
    .ZN(_06712_));
 NOR2_X1 _23849_ (.A1(net375),
    .A2(_06390_),
    .ZN(_06713_));
 AOI21_X2 _23850_ (.A(_06713_),
    .B1(_06399_),
    .B2(_03824_),
    .ZN(_06714_));
 OAI211_X2 _23851_ (.A(_03404_),
    .B(_06712_),
    .C1(_06714_),
    .C2(_06378_),
    .ZN(_06715_));
 AOI22_X1 _23852_ (.A1(_13259_),
    .A2(_06379_),
    .B1(_06710_),
    .B2(_06715_),
    .ZN(_06716_));
 MUX2_X1 _23853_ (.A(_04811_),
    .B(_06716_),
    .S(_03440_),
    .Z(_06717_));
 MUX2_X1 _23854_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B(_06717_),
    .S(_06383_),
    .Z(_01331_));
 NAND3_X1 _23855_ (.A1(_03450_),
    .A2(_05089_),
    .A3(_06383_),
    .ZN(_06718_));
 AOI221_X2 _23856_ (.A(_06452_),
    .B1(_06714_),
    .B2(_03403_),
    .C1(_03650_),
    .C2(\alu_adder_result_ex[28] ),
    .ZN(_06719_));
 AOI21_X1 _23857_ (.A(_06719_),
    .B1(_06379_),
    .B2(_03131_),
    .ZN(_06720_));
 NOR2_X1 _23858_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_06391_),
    .ZN(_06721_));
 AOI21_X2 _23859_ (.A(_06721_),
    .B1(_06473_),
    .B2(_03827_),
    .ZN(_06722_));
 NOR2_X1 _23860_ (.A1(_06378_),
    .A2(_06722_),
    .ZN(_06723_));
 INV_X1 _23861_ (.A(_00096_),
    .ZN(_06724_));
 INV_X1 _23862_ (.A(_06570_),
    .ZN(_06725_));
 AOI21_X2 _23863_ (.A(_06724_),
    .B1(_06725_),
    .B2(_06614_),
    .ZN(_06726_));
 AOI21_X1 _23864_ (.A(_06723_),
    .B1(_06726_),
    .B2(_06387_),
    .ZN(_06727_));
 AOI21_X1 _23865_ (.A(_06720_),
    .B1(_06727_),
    .B2(_06385_),
    .ZN(_06728_));
 INV_X1 _23866_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .ZN(_06729_));
 OAI221_X1 _23867_ (.A(_06718_),
    .B1(_06728_),
    .B2(_06670_),
    .C1(_06729_),
    .C2(_06383_),
    .ZN(_01332_));
 AOI22_X1 _23868_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(_06450_),
    .B1(_06598_),
    .B2(_05111_),
    .ZN(_06730_));
 AOI221_X2 _23869_ (.A(_06453_),
    .B1(_06722_),
    .B2(_03431_),
    .C1(_03651_),
    .C2(net14),
    .ZN(_06731_));
 INV_X1 _23870_ (.A(_06731_),
    .ZN(_06732_));
 OAI21_X1 _23871_ (.A(_00097_),
    .B1(_06570_),
    .B2(_06621_),
    .ZN(_06733_));
 MUX2_X1 _23872_ (.A(net14),
    .B(_03829_),
    .S(_06399_),
    .Z(_06734_));
 MUX2_X1 _23873_ (.A(_06733_),
    .B(_06734_),
    .S(_06396_),
    .Z(_06735_));
 AOI21_X1 _23874_ (.A(_06732_),
    .B1(_06735_),
    .B2(_06385_),
    .ZN(_06736_));
 OAI21_X1 _23875_ (.A(_06375_),
    .B1(_06564_),
    .B2(_03769_),
    .ZN(_06737_));
 OAI21_X1 _23876_ (.A(_06730_),
    .B1(_06736_),
    .B2(_06737_),
    .ZN(_01333_));
 NAND2_X1 _23877_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_06450_),
    .ZN(_06738_));
 AOI221_X1 _23878_ (.A(_06453_),
    .B1(_06734_),
    .B2(_03403_),
    .C1(_03650_),
    .C2(\alu_adder_result_ex[30] ),
    .ZN(_06739_));
 INV_X1 _23879_ (.A(_06739_),
    .ZN(_06740_));
 OAI21_X1 _23880_ (.A(_00098_),
    .B1(_06570_),
    .B2(_06630_),
    .ZN(_06741_));
 MUX2_X1 _23881_ (.A(\alu_adder_result_ex[30] ),
    .B(_03831_),
    .S(_06473_),
    .Z(_06742_));
 MUX2_X1 _23882_ (.A(_06741_),
    .B(_06742_),
    .S(_06396_),
    .Z(_06743_));
 AOI21_X1 _23883_ (.A(_06740_),
    .B1(_06743_),
    .B2(_06385_),
    .ZN(_06744_));
 OAI21_X1 _23884_ (.A(_03440_),
    .B1(_06564_),
    .B2(_03311_),
    .ZN(_06745_));
 OR2_X1 _23885_ (.A1(_06374_),
    .A2(_06745_),
    .ZN(_06746_));
 OAI221_X1 _23886_ (.A(_06738_),
    .B1(_06744_),
    .B2(_06746_),
    .C1(_06671_),
    .C2(_05173_),
    .ZN(_01334_));
 NAND2_X1 _23887_ (.A1(_04791_),
    .A2(_05223_),
    .ZN(_06747_));
 OAI21_X1 _23888_ (.A(_06747_),
    .B1(_05219_),
    .B2(_04791_),
    .ZN(_06748_));
 AOI22_X1 _23889_ (.A1(_03408_),
    .A2(_06450_),
    .B1(_06598_),
    .B2(_06748_),
    .ZN(_06749_));
 OAI21_X2 _23890_ (.A(_06366_),
    .B1(_03417_),
    .B2(_04044_),
    .ZN(_06750_));
 OAI21_X1 _23891_ (.A(_00099_),
    .B1(_06570_),
    .B2(_06639_),
    .ZN(_06751_));
 AND2_X1 _23892_ (.A1(_03408_),
    .A2(net279),
    .ZN(_06752_));
 MUX2_X1 _23893_ (.A(_06751_),
    .B(_06752_),
    .S(_06395_),
    .Z(_06753_));
 AOI221_X2 _23894_ (.A(_06750_),
    .B1(_06753_),
    .B2(_03404_),
    .C1(_06742_),
    .C2(_03614_),
    .ZN(_06754_));
 OAI21_X1 _23895_ (.A(_06375_),
    .B1(_06564_),
    .B2(_03783_),
    .ZN(_06755_));
 OAI21_X1 _23896_ (.A(_06749_),
    .B1(_06754_),
    .B2(_06755_),
    .ZN(_01335_));
 INV_X1 _23897_ (.A(_15822_),
    .ZN(_06756_));
 NAND3_X1 _23898_ (.A1(_15811_),
    .A2(_05107_),
    .A3(_05161_),
    .ZN(_06757_));
 AOI21_X1 _23899_ (.A(_05170_),
    .B1(_05166_),
    .B2(_06757_),
    .ZN(_06758_));
 OAI21_X1 _23900_ (.A(_15823_),
    .B1(_15816_),
    .B2(_06758_),
    .ZN(_06759_));
 AND2_X1 _23901_ (.A1(_06756_),
    .A2(_06759_),
    .ZN(_06760_));
 XNOR2_X1 _23902_ (.A(_15830_),
    .B(_06760_),
    .ZN(_06761_));
 NAND3_X1 _23903_ (.A1(_03450_),
    .A2(_04791_),
    .A3(_06761_),
    .ZN(_06762_));
 AOI22_X2 _23904_ (.A1(_06453_),
    .A2(_06378_),
    .B1(_06752_),
    .B2(_03614_),
    .ZN(_06763_));
 OAI21_X1 _23905_ (.A(_06762_),
    .B1(_06763_),
    .B2(_03450_),
    .ZN(_06764_));
 MUX2_X1 _23906_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B(_06764_),
    .S(_06383_),
    .Z(_01336_));
 AOI21_X1 _23907_ (.A(_06450_),
    .B1(_06387_),
    .B2(_06453_),
    .ZN(_06765_));
 NOR2_X1 _23908_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A2(_06383_),
    .ZN(_06766_));
 NAND4_X1 _23909_ (.A1(_10888_),
    .A2(_03450_),
    .A3(_04791_),
    .A4(_06383_),
    .ZN(_06767_));
 XOR2_X1 _23910_ (.A(_15344_),
    .B(_15732_),
    .Z(_06768_));
 XNOR2_X1 _23911_ (.A(_15340_),
    .B(_06768_),
    .ZN(_06769_));
 XOR2_X1 _23912_ (.A(_15347_),
    .B(_14815_),
    .Z(_06770_));
 XNOR2_X1 _23913_ (.A(_15335_),
    .B(_15826_),
    .ZN(_06771_));
 XNOR2_X1 _23914_ (.A(_06770_),
    .B(_06771_),
    .ZN(_06772_));
 XNOR2_X1 _23915_ (.A(_15261_),
    .B(_15304_),
    .ZN(_06773_));
 XNOR2_X1 _23916_ (.A(_06772_),
    .B(_06773_),
    .ZN(_06774_));
 XOR2_X1 _23917_ (.A(_15327_),
    .B(_15220_),
    .Z(_06775_));
 XNOR2_X1 _23918_ (.A(_15326_),
    .B(_15350_),
    .ZN(_06776_));
 XNOR2_X1 _23919_ (.A(_06775_),
    .B(_06776_),
    .ZN(_06777_));
 XNOR2_X1 _23920_ (.A(_15332_),
    .B(_15338_),
    .ZN(_06778_));
 XNOR2_X1 _23921_ (.A(_15303_),
    .B(_15330_),
    .ZN(_06779_));
 XNOR2_X1 _23922_ (.A(_06778_),
    .B(_06779_),
    .ZN(_06780_));
 XNOR2_X1 _23923_ (.A(_06777_),
    .B(_06780_),
    .ZN(_06781_));
 XNOR2_X1 _23924_ (.A(_06774_),
    .B(_06781_),
    .ZN(_06782_));
 XNOR2_X1 _23925_ (.A(_06769_),
    .B(_06782_),
    .ZN(_06783_));
 OAI21_X1 _23926_ (.A(_03802_),
    .B1(_03794_),
    .B2(_00132_),
    .ZN(_06784_));
 NAND2_X1 _23927_ (.A1(_03664_),
    .A2(_06784_),
    .ZN(_06785_));
 XNOR2_X1 _23928_ (.A(_06783_),
    .B(_06785_),
    .ZN(_06786_));
 INV_X1 _23929_ (.A(_15823_),
    .ZN(_06787_));
 OAI21_X1 _23930_ (.A(_06756_),
    .B1(_05222_),
    .B2(_06787_),
    .ZN(_06788_));
 AOI21_X1 _23931_ (.A(_15829_),
    .B1(_06788_),
    .B2(_15830_),
    .ZN(_06789_));
 XNOR2_X1 _23932_ (.A(_06786_),
    .B(_06789_),
    .ZN(_06790_));
 OAI22_X1 _23933_ (.A1(_06765_),
    .A2(_06766_),
    .B1(_06767_),
    .B2(_06790_),
    .ZN(_01337_));
 MUX2_X1 _23934_ (.A(\alu_adder_result_ex[6] ),
    .B(_11158_),
    .S(_03779_),
    .Z(_06791_));
 MUX2_X1 _23935_ (.A(_06791_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .S(_03612_),
    .Z(_01338_));
 MUX2_X1 _23936_ (.A(\alu_adder_result_ex[7] ),
    .B(_11202_),
    .S(_03779_),
    .Z(_06792_));
 MUX2_X1 _23937_ (.A(_06792_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .S(_03612_),
    .Z(_01339_));
 NAND2_X1 _23938_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .A2(_03613_),
    .ZN(_06793_));
 NAND2_X1 _23939_ (.A1(_11241_),
    .A2(_03780_),
    .ZN(_06794_));
 OAI21_X1 _23940_ (.A(_06794_),
    .B1(_03780_),
    .B2(\alu_adder_result_ex[8] ),
    .ZN(_06795_));
 OAI21_X1 _23941_ (.A(_06793_),
    .B1(_06795_),
    .B2(_03613_),
    .ZN(_01340_));
 MUX2_X1 _23942_ (.A(\alu_adder_result_ex[9] ),
    .B(_03727_),
    .S(_03779_),
    .Z(_06796_));
 MUX2_X1 _23943_ (.A(_06796_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .S(_03612_),
    .Z(_01341_));
 NOR2_X4 _23944_ (.A1(_03836_),
    .A2(_03921_),
    .ZN(_06797_));
 NAND2_X1 _23945_ (.A1(\cs_registers_i.csr_mepc_o[4] ),
    .A2(_06797_),
    .ZN(_06798_));
 NAND2_X2 _23946_ (.A1(_03918_),
    .A2(_03867_),
    .ZN(_06799_));
 NAND3_X1 _23947_ (.A1(_03863_),
    .A2(_03864_),
    .A3(_06799_),
    .ZN(_06800_));
 NAND2_X1 _23948_ (.A1(_03856_),
    .A2(_03857_),
    .ZN(_06801_));
 AOI221_X2 _23949_ (.A(_06800_),
    .B1(_03866_),
    .B2(_03902_),
    .C1(_06801_),
    .C2(_03900_),
    .ZN(_06802_));
 OR3_X4 _23950_ (.A1(_03465_),
    .A2(_03839_),
    .A3(_03921_),
    .ZN(_06803_));
 OAI221_X2 _23951_ (.A(_06798_),
    .B1(_06802_),
    .B2(_03873_),
    .C1(_01164_),
    .C2(_06803_),
    .ZN(_06804_));
 OR2_X1 _23952_ (.A1(_03889_),
    .A2(_06804_),
    .ZN(_06805_));
 AOI21_X4 _23953_ (.A(_06805_),
    .B1(\alu_adder_result_ex[4] ),
    .B2(_03929_),
    .ZN(_06806_));
 NOR2_X2 _23954_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .A2(_03936_),
    .ZN(_06807_));
 NOR2_X2 _23955_ (.A1(_06806_),
    .A2(_06807_),
    .ZN(_06808_));
 NAND3_X1 _23956_ (.A1(net135),
    .A2(\cs_registers_i.mie_q[15] ),
    .A3(_03860_),
    .ZN(_06809_));
 AND2_X1 _23957_ (.A1(_03865_),
    .A2(_06799_),
    .ZN(_06810_));
 AOI21_X2 _23958_ (.A(_03873_),
    .B1(_06809_),
    .B2(_06810_),
    .ZN(_06811_));
 INV_X1 _23959_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .ZN(_06812_));
 OAI22_X2 _23960_ (.A1(_06812_),
    .A2(_03894_),
    .B1(_03895_),
    .B2(_01165_),
    .ZN(_06813_));
 NOR2_X1 _23961_ (.A1(_03952_),
    .A2(_03891_),
    .ZN(_06814_));
 AOI221_X2 _23962_ (.A(_06811_),
    .B1(_06813_),
    .B2(_06814_),
    .C1(\alu_adder_result_ex[5] ),
    .C2(net22),
    .ZN(_06815_));
 AND2_X2 _23963_ (.A1(_03935_),
    .A2(_06815_),
    .ZN(_06816_));
 INV_X1 _23964_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .ZN(_06817_));
 AOI21_X4 _23965_ (.A(_06816_),
    .B1(_03957_),
    .B2(_06817_),
    .ZN(_06818_));
 NAND3_X2 _23966_ (.A1(_16111_),
    .A2(_06808_),
    .A3(_06818_),
    .ZN(_06819_));
 OAI21_X2 _23967_ (.A(_03436_),
    .B1(_03954_),
    .B2(_03838_),
    .ZN(_06820_));
 NAND2_X4 _23968_ (.A1(_03459_),
    .A2(_06820_),
    .ZN(_06821_));
 NOR2_X1 _23969_ (.A1(_01167_),
    .A2(_06821_),
    .ZN(_06822_));
 AOI221_X2 _23970_ (.A(_06822_),
    .B1(_03922_),
    .B2(\cs_registers_i.csr_mepc_o[8] ),
    .C1(\cs_registers_i.csr_depc_o[8] ),
    .C2(_03925_),
    .ZN(_06823_));
 NAND2_X1 _23971_ (.A1(net34),
    .A2(_03897_),
    .ZN(_06824_));
 NAND3_X2 _23972_ (.A1(_03935_),
    .A2(_06823_),
    .A3(_06824_),
    .ZN(_06825_));
 AOI21_X4 _23973_ (.A(_06825_),
    .B1(\alu_adder_result_ex[8] ),
    .B2(_03929_),
    .ZN(_06826_));
 INV_X1 _23974_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .ZN(_06827_));
 AOI21_X4 _23975_ (.A(_06826_),
    .B1(_03957_),
    .B2(_06827_),
    .ZN(_06828_));
 NOR2_X1 _23976_ (.A1(_01168_),
    .A2(_06821_),
    .ZN(_06829_));
 AOI221_X2 _23977_ (.A(_06829_),
    .B1(_03922_),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .C1(\cs_registers_i.csr_depc_o[9] ),
    .C2(_03925_),
    .ZN(_06830_));
 NAND2_X1 _23978_ (.A1(net22),
    .A2(\alu_adder_result_ex[9] ),
    .ZN(_06831_));
 NAND2_X1 _23979_ (.A1(_06830_),
    .A2(_06831_),
    .ZN(_06832_));
 NOR2_X1 _23980_ (.A1(net22),
    .A2(_03893_),
    .ZN(_06833_));
 NAND2_X2 _23981_ (.A1(_03461_),
    .A2(_03896_),
    .ZN(_06834_));
 NAND2_X4 _23982_ (.A1(_06833_),
    .A2(_06834_),
    .ZN(_06835_));
 MUX2_X1 _23983_ (.A(net35),
    .B(_06832_),
    .S(_06835_),
    .Z(_06836_));
 NAND2_X1 _23984_ (.A1(_03936_),
    .A2(_06836_),
    .ZN(_06837_));
 INV_X1 _23985_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .ZN(_06838_));
 OAI21_X2 _23986_ (.A(_06837_),
    .B1(_03936_),
    .B2(_06838_),
    .ZN(_06839_));
 NOR2_X2 _23987_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .A2(_03935_),
    .ZN(_06840_));
 NAND2_X1 _23988_ (.A1(net22),
    .A2(\alu_adder_result_ex[7] ),
    .ZN(_06841_));
 AOI22_X2 _23989_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_03922_),
    .B1(_03925_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .ZN(_06842_));
 AND3_X2 _23990_ (.A1(_03898_),
    .A2(_06841_),
    .A3(_06842_),
    .ZN(_06843_));
 AOI21_X4 _23991_ (.A(_03873_),
    .B1(_06799_),
    .B2(_03902_),
    .ZN(_06844_));
 AOI221_X2 _23992_ (.A(_06844_),
    .B1(_03922_),
    .B2(\cs_registers_i.csr_mepc_o[6] ),
    .C1(_05601_),
    .C2(_03925_),
    .ZN(_06845_));
 NAND2_X1 _23993_ (.A1(_03935_),
    .A2(_06845_),
    .ZN(_06846_));
 AOI21_X4 _23994_ (.A(_06846_),
    .B1(\alu_adder_result_ex[6] ),
    .B2(_03929_),
    .ZN(_06847_));
 NOR2_X2 _23995_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(_03935_),
    .ZN(_06848_));
 NOR4_X4 _23996_ (.A1(_06840_),
    .A2(_06843_),
    .A3(_06847_),
    .A4(_06848_),
    .ZN(_06849_));
 NAND3_X1 _23997_ (.A1(_06828_),
    .A2(_06839_),
    .A3(_06849_),
    .ZN(_06850_));
 OR2_X1 _23998_ (.A1(_06819_),
    .A2(_06850_),
    .ZN(_06851_));
 BUF_X4 _23999_ (.A(_04154_),
    .Z(_06852_));
 AOI22_X1 _24000_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(_03922_),
    .B1(_03925_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .ZN(_06853_));
 OAI21_X1 _24001_ (.A(_06853_),
    .B1(_06821_),
    .B2(_01169_),
    .ZN(_06854_));
 AOI221_X2 _24002_ (.A(_06854_),
    .B1(\alu_adder_result_ex[10] ),
    .B2(_03929_),
    .C1(net3),
    .C2(_03897_),
    .ZN(_06855_));
 OR2_X1 _24003_ (.A1(_06852_),
    .A2(_06855_),
    .ZN(_06856_));
 XOR2_X1 _24004_ (.A(_06851_),
    .B(_06856_),
    .Z(_06857_));
 BUF_X4 _24005_ (.A(_06852_),
    .Z(_06858_));
 AOI21_X1 _24006_ (.A(_06857_),
    .B1(_06858_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .ZN(_06859_));
 INV_X1 _24007_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .ZN(_06860_));
 OR3_X1 _24008_ (.A1(_06860_),
    .A2(_04164_),
    .A3(_06851_),
    .ZN(_06861_));
 OAI21_X1 _24009_ (.A(_06861_),
    .B1(_16107_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .ZN(_06862_));
 CLKBUF_X3 _24010_ (.A(_06858_),
    .Z(_06863_));
 AOI21_X1 _24011_ (.A(_06859_),
    .B1(_06862_),
    .B2(_06863_),
    .ZN(_01342_));
 NAND3_X1 _24012_ (.A1(_00550_),
    .A2(_03844_),
    .A3(_03953_),
    .ZN(_06864_));
 OR3_X1 _24013_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_03878_),
    .A3(_03953_),
    .ZN(_06865_));
 NAND3_X1 _24014_ (.A1(_03893_),
    .A2(_06864_),
    .A3(_06865_),
    .ZN(_06866_));
 AOI22_X1 _24015_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_03922_),
    .B1(_03925_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .ZN(_06867_));
 NAND2_X1 _24016_ (.A1(_06866_),
    .A2(_06867_),
    .ZN(_06868_));
 AOI221_X2 _24017_ (.A(_06868_),
    .B1(\alu_adder_result_ex[11] ),
    .B2(net22),
    .C1(net4),
    .C2(_03897_),
    .ZN(_06869_));
 NOR2_X1 _24018_ (.A1(_03957_),
    .A2(_06869_),
    .ZN(_06870_));
 AOI21_X2 _24019_ (.A(_06870_),
    .B1(_03957_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .ZN(_06871_));
 MUX2_X2 _24020_ (.A(_06860_),
    .B(_06855_),
    .S(_03936_),
    .Z(_06872_));
 INV_X1 _24021_ (.A(_16109_),
    .ZN(_06873_));
 NAND2_X1 _24022_ (.A1(_16110_),
    .A2(_06818_),
    .ZN(_06874_));
 NOR4_X4 _24023_ (.A1(_06873_),
    .A2(_06806_),
    .A3(_06807_),
    .A4(_06874_),
    .ZN(_06875_));
 NAND4_X1 _24024_ (.A1(_06828_),
    .A2(_06839_),
    .A3(_06849_),
    .A4(_06875_),
    .ZN(_06876_));
 NOR2_X1 _24025_ (.A1(_06872_),
    .A2(_06876_),
    .ZN(_06877_));
 XNOR2_X1 _24026_ (.A(_06871_),
    .B(_06877_),
    .ZN(_06878_));
 NAND2_X2 _24027_ (.A1(_06852_),
    .A2(_04164_),
    .ZN(_06879_));
 CLKBUF_X3 _24028_ (.A(_06879_),
    .Z(_06880_));
 MUX2_X1 _24029_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .B(_06878_),
    .S(_06880_),
    .Z(_01343_));
 INV_X1 _24030_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .ZN(_06881_));
 OR4_X2 _24031_ (.A1(_06819_),
    .A2(_06850_),
    .A3(_06871_),
    .A4(_06872_),
    .ZN(_06882_));
 NOR2_X1 _24032_ (.A1(_04164_),
    .A2(_06882_),
    .ZN(_06883_));
 XNOR2_X1 _24033_ (.A(_06881_),
    .B(_06883_),
    .ZN(_06884_));
 NAND2_X1 _24034_ (.A1(_03931_),
    .A2(\alu_adder_result_ex[12] ),
    .ZN(_06885_));
 AOI22_X2 _24035_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(_03922_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .ZN(_06886_));
 OAI21_X2 _24036_ (.A(_06886_),
    .B1(_06821_),
    .B2(_00549_),
    .ZN(_06887_));
 BUF_X4 _24037_ (.A(_03897_),
    .Z(_06888_));
 BUF_X4 _24038_ (.A(_06888_),
    .Z(_06889_));
 AOI21_X1 _24039_ (.A(_06887_),
    .B1(_06889_),
    .B2(net5),
    .ZN(_06890_));
 NAND2_X1 _24040_ (.A1(_06885_),
    .A2(_06890_),
    .ZN(_06891_));
 XNOR2_X1 _24041_ (.A(_06882_),
    .B(_06891_),
    .ZN(_06892_));
 BUF_X4 _24042_ (.A(_03939_),
    .Z(_06893_));
 MUX2_X1 _24043_ (.A(_06884_),
    .B(_06892_),
    .S(_06893_),
    .Z(_01344_));
 AOI22_X1 _24044_ (.A1(\cs_registers_i.csr_mepc_o[13] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[13] ),
    .ZN(_06894_));
 BUF_X4 _24045_ (.A(_06821_),
    .Z(_06895_));
 OAI21_X1 _24046_ (.A(_06894_),
    .B1(_06895_),
    .B2(_01170_),
    .ZN(_06896_));
 AOI21_X2 _24047_ (.A(_06896_),
    .B1(_06888_),
    .B2(net6),
    .ZN(_06897_));
 NAND2_X1 _24048_ (.A1(_03936_),
    .A2(_06897_),
    .ZN(_06898_));
 AOI21_X2 _24049_ (.A(_06898_),
    .B1(\alu_adder_result_ex[13] ),
    .B2(_03930_),
    .ZN(_06899_));
 INV_X1 _24050_ (.A(_06899_),
    .ZN(_06900_));
 OAI21_X2 _24051_ (.A(_06900_),
    .B1(_03938_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .ZN(_06901_));
 NAND2_X1 _24052_ (.A1(_06828_),
    .A2(_06849_),
    .ZN(_06902_));
 AOI221_X2 _24053_ (.A(_06887_),
    .B1(\alu_adder_result_ex[12] ),
    .B2(_03929_),
    .C1(net5),
    .C2(_06888_),
    .ZN(_06903_));
 MUX2_X2 _24054_ (.A(_06881_),
    .B(_06903_),
    .S(_03937_),
    .Z(_06904_));
 OR2_X1 _24055_ (.A1(_04154_),
    .A2(_06869_),
    .ZN(_06905_));
 INV_X1 _24056_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .ZN(_06906_));
 OAI21_X1 _24057_ (.A(_06905_),
    .B1(_03937_),
    .B2(_06906_),
    .ZN(_06907_));
 NAND3_X1 _24058_ (.A1(_06839_),
    .A2(_06907_),
    .A3(_06875_),
    .ZN(_06908_));
 NOR4_X4 _24059_ (.A1(_06902_),
    .A2(_06872_),
    .A3(_06904_),
    .A4(_06908_),
    .ZN(_06909_));
 XNOR2_X1 _24060_ (.A(_06901_),
    .B(_06909_),
    .ZN(_06910_));
 MUX2_X1 _24061_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .B(_06910_),
    .S(_06880_),
    .Z(_01345_));
 NOR3_X4 _24062_ (.A1(_06882_),
    .A2(_06901_),
    .A3(_06904_),
    .ZN(_06911_));
 NAND3_X1 _24063_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(_16107_),
    .A3(_06911_),
    .ZN(_06912_));
 OAI21_X1 _24064_ (.A(_06912_),
    .B1(_16107_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .ZN(_06913_));
 NAND2_X1 _24065_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(_04154_),
    .ZN(_06914_));
 AOI22_X1 _24066_ (.A1(\cs_registers_i.csr_mepc_o[14] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[14] ),
    .ZN(_06915_));
 OAI21_X1 _24067_ (.A(_06915_),
    .B1(_06895_),
    .B2(_01171_),
    .ZN(_06916_));
 AOI221_X2 _24068_ (.A(_06916_),
    .B1(\alu_adder_result_ex[14] ),
    .B2(_03929_),
    .C1(net7),
    .C2(_06888_),
    .ZN(_06917_));
 OR2_X4 _24069_ (.A1(_04154_),
    .A2(_06917_),
    .ZN(_06918_));
 XOR2_X1 _24070_ (.A(_06911_),
    .B(_06918_),
    .Z(_06919_));
 AOI22_X1 _24071_ (.A1(_06863_),
    .A2(_06913_),
    .B1(_06914_),
    .B2(_06919_),
    .ZN(_01346_));
 NOR3_X4 _24072_ (.A1(_11426_),
    .A2(_12266_),
    .A3(_12273_),
    .ZN(_06920_));
 AOI22_X1 _24073_ (.A1(\cs_registers_i.csr_mepc_o[15] ),
    .A2(_03469_),
    .B1(_03476_),
    .B2(\cs_registers_i.csr_depc_o[15] ),
    .ZN(_06921_));
 OAI22_X1 _24074_ (.A1(_01172_),
    .A2(_06821_),
    .B1(_06921_),
    .B2(_03921_),
    .ZN(_06922_));
 OR3_X1 _24075_ (.A1(_06888_),
    .A2(_06920_),
    .A3(_06922_),
    .ZN(_06923_));
 OAI221_X2 _24076_ (.A(_06923_),
    .B1(_03888_),
    .B2(_03883_),
    .C1(net8),
    .C2(_06835_),
    .ZN(_06924_));
 INV_X1 _24077_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .ZN(_06925_));
 OAI21_X2 _24078_ (.A(_06924_),
    .B1(_03936_),
    .B2(_06925_),
    .ZN(_06926_));
 INV_X1 _24079_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .ZN(_06927_));
 AOI21_X2 _24080_ (.A(_06899_),
    .B1(_06852_),
    .B2(_06927_),
    .ZN(_06928_));
 NAND2_X4 _24081_ (.A1(_06914_),
    .A2(_06918_),
    .ZN(_06929_));
 NAND3_X2 _24082_ (.A1(_06928_),
    .A2(_06909_),
    .A3(_06929_),
    .ZN(_06930_));
 XNOR2_X1 _24083_ (.A(_06926_),
    .B(_06930_),
    .ZN(_06931_));
 MUX2_X1 _24084_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .B(_06931_),
    .S(_06880_),
    .Z(_01347_));
 NOR2_X1 _24085_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A2(_03936_),
    .ZN(_06932_));
 NAND3_X1 _24086_ (.A1(_03844_),
    .A2(_01173_),
    .A3(_03953_),
    .ZN(_06933_));
 OR3_X1 _24087_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_03878_),
    .A3(_03953_),
    .ZN(_06934_));
 NAND3_X1 _24088_ (.A1(_03893_),
    .A2(_06933_),
    .A3(_06934_),
    .ZN(_06935_));
 AOI22_X1 _24089_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .ZN(_06936_));
 NAND2_X1 _24090_ (.A1(net9),
    .A2(_06888_),
    .ZN(_06937_));
 AND4_X2 _24091_ (.A1(_03936_),
    .A2(_06935_),
    .A3(_06936_),
    .A4(_06937_),
    .ZN(_06938_));
 NAND3_X2 _24092_ (.A1(_03930_),
    .A2(_12445_),
    .A3(_12446_),
    .ZN(_06939_));
 AOI21_X4 _24093_ (.A(_06932_),
    .B1(_06938_),
    .B2(_06939_),
    .ZN(_06940_));
 AND3_X1 _24094_ (.A1(_06911_),
    .A2(_06929_),
    .A3(_06926_),
    .ZN(_06941_));
 XOR2_X1 _24095_ (.A(_06940_),
    .B(_06941_),
    .Z(_06942_));
 MUX2_X1 _24096_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .B(_06942_),
    .S(_06880_),
    .Z(_01348_));
 NAND2_X1 _24097_ (.A1(_06926_),
    .A2(_06940_),
    .ZN(_06943_));
 NOR2_X1 _24098_ (.A1(_06930_),
    .A2(_06943_),
    .ZN(_06944_));
 NAND2_X1 _24099_ (.A1(_16107_),
    .A2(_06944_),
    .ZN(_06945_));
 XNOR2_X1 _24100_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .B(_06945_),
    .ZN(_06946_));
 AOI22_X2 _24101_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(_03469_),
    .B1(_03476_),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .ZN(_06947_));
 OAI22_X2 _24102_ (.A1(_01174_),
    .A2(_06821_),
    .B1(_06947_),
    .B2(_03921_),
    .ZN(_06948_));
 AOI21_X1 _24103_ (.A(_06948_),
    .B1(\alu_adder_result_ex[17] ),
    .B2(_03929_),
    .ZN(_06949_));
 NAND2_X1 _24104_ (.A1(_06835_),
    .A2(_06949_),
    .ZN(_06950_));
 OAI21_X2 _24105_ (.A(_06950_),
    .B1(_06835_),
    .B2(net10),
    .ZN(_06951_));
 XNOR2_X1 _24106_ (.A(_06944_),
    .B(_06951_),
    .ZN(_06952_));
 MUX2_X1 _24107_ (.A(_06946_),
    .B(_06952_),
    .S(_06893_),
    .Z(_01349_));
 NOR2_X1 _24108_ (.A1(net11),
    .A2(_06835_),
    .ZN(_06953_));
 INV_X1 _24109_ (.A(\cs_registers_i.csr_depc_o[18] ),
    .ZN(_06954_));
 OAI22_X2 _24110_ (.A1(_06954_),
    .A2(_06803_),
    .B1(_06895_),
    .B2(_01175_),
    .ZN(_06955_));
 AOI21_X2 _24111_ (.A(_06955_),
    .B1(_06797_),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .ZN(_06956_));
 NAND2_X1 _24112_ (.A1(_06835_),
    .A2(_06956_),
    .ZN(_06957_));
 AOI21_X2 _24113_ (.A(_06957_),
    .B1(\alu_adder_result_ex[18] ),
    .B2(_03930_),
    .ZN(_06958_));
 OR3_X1 _24114_ (.A1(_06852_),
    .A2(_06953_),
    .A3(_06958_),
    .ZN(_06959_));
 INV_X1 _24115_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .ZN(_06960_));
 OAI21_X2 _24116_ (.A(_06959_),
    .B1(_03938_),
    .B2(_06960_),
    .ZN(_06961_));
 NAND2_X1 _24117_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(_03957_),
    .ZN(_06962_));
 OAI21_X1 _24118_ (.A(_06962_),
    .B1(_06951_),
    .B2(_04154_),
    .ZN(_06963_));
 AND3_X1 _24119_ (.A1(_06926_),
    .A2(_06940_),
    .A3(_06963_),
    .ZN(_06964_));
 AND3_X1 _24120_ (.A1(_06911_),
    .A2(_06929_),
    .A3(_06964_),
    .ZN(_06965_));
 XOR2_X1 _24121_ (.A(_06961_),
    .B(_06965_),
    .Z(_06966_));
 MUX2_X1 _24122_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .B(_06966_),
    .S(_06880_),
    .Z(_01350_));
 AND2_X1 _24123_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(_03957_),
    .ZN(_06967_));
 NOR4_X1 _24124_ (.A1(_06871_),
    .A2(_06872_),
    .A3(_06876_),
    .A4(_06904_),
    .ZN(_06968_));
 AND3_X1 _24125_ (.A1(_06928_),
    .A2(_06968_),
    .A3(_06929_),
    .ZN(_06969_));
 NAND3_X1 _24126_ (.A1(_06969_),
    .A2(_06961_),
    .A3(_06964_),
    .ZN(_06970_));
 OAI21_X1 _24127_ (.A(_06967_),
    .B1(_06970_),
    .B2(_04164_),
    .ZN(_06971_));
 AOI22_X1 _24128_ (.A1(\cs_registers_i.csr_mepc_o[19] ),
    .A2(_03922_),
    .B1(_03925_),
    .B2(\cs_registers_i.csr_depc_o[19] ),
    .ZN(_06972_));
 OAI21_X1 _24129_ (.A(_06972_),
    .B1(_06821_),
    .B2(_01176_),
    .ZN(_06973_));
 AOI221_X2 _24130_ (.A(_06973_),
    .B1(\alu_adder_result_ex[19] ),
    .B2(_03929_),
    .C1(net12),
    .C2(_06888_),
    .ZN(_06974_));
 NOR2_X2 _24131_ (.A1(_03957_),
    .A2(_06974_),
    .ZN(_06975_));
 INV_X1 _24132_ (.A(_06975_),
    .ZN(_06976_));
 NAND2_X1 _24133_ (.A1(_06970_),
    .A2(_06976_),
    .ZN(_06977_));
 NAND2_X1 _24134_ (.A1(_06880_),
    .A2(_06977_),
    .ZN(_06978_));
 INV_X1 _24135_ (.A(_06967_),
    .ZN(_06979_));
 AOI21_X1 _24136_ (.A(_06970_),
    .B1(_06976_),
    .B2(_06979_),
    .ZN(_06980_));
 OAI21_X1 _24137_ (.A(_06971_),
    .B1(_06978_),
    .B2(_06980_),
    .ZN(_01351_));
 INV_X1 _24138_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .ZN(_06981_));
 OAI21_X1 _24139_ (.A(_06975_),
    .B1(_06835_),
    .B2(net11),
    .ZN(_06982_));
 OAI22_X2 _24140_ (.A1(_06960_),
    .A2(_06979_),
    .B1(_06982_),
    .B2(_06958_),
    .ZN(_06983_));
 AND2_X1 _24141_ (.A1(_06964_),
    .A2(_06983_),
    .ZN(_06984_));
 NAND3_X1 _24142_ (.A1(_06911_),
    .A2(_06929_),
    .A3(_06984_),
    .ZN(_06985_));
 NOR2_X1 _24143_ (.A1(_04164_),
    .A2(_06985_),
    .ZN(_06986_));
 XNOR2_X1 _24144_ (.A(_06981_),
    .B(_06986_),
    .ZN(_06987_));
 NOR4_X4 _24145_ (.A1(_11426_),
    .A2(_12776_),
    .A3(_12778_),
    .A4(_12781_),
    .ZN(_06988_));
 BUF_X4 _24146_ (.A(_03953_),
    .Z(_06989_));
 NAND3_X1 _24147_ (.A1(_03844_),
    .A2(_01177_),
    .A3(_06989_),
    .ZN(_06990_));
 OR3_X1 _24148_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_03878_),
    .A3(_03953_),
    .ZN(_06991_));
 NAND3_X1 _24149_ (.A1(_03893_),
    .A2(_06990_),
    .A3(_06991_),
    .ZN(_06992_));
 AOI22_X2 _24150_ (.A1(\cs_registers_i.csr_mepc_o[20] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .ZN(_06993_));
 NAND2_X1 _24151_ (.A1(net13),
    .A2(_06888_),
    .ZN(_06994_));
 NAND3_X2 _24152_ (.A1(_06992_),
    .A2(_06993_),
    .A3(_06994_),
    .ZN(_06995_));
 NOR2_X1 _24153_ (.A1(_06988_),
    .A2(_06995_),
    .ZN(_06996_));
 XOR2_X1 _24154_ (.A(_06985_),
    .B(_06996_),
    .Z(_06997_));
 BUF_X4 _24155_ (.A(_03939_),
    .Z(_06998_));
 MUX2_X1 _24156_ (.A(_06987_),
    .B(_06997_),
    .S(_06998_),
    .Z(_01352_));
 NOR2_X1 _24157_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .A2(_06880_),
    .ZN(_06999_));
 INV_X1 _24158_ (.A(\cs_registers_i.csr_depc_o[21] ),
    .ZN(_07000_));
 OAI22_X2 _24159_ (.A1(_07000_),
    .A2(_06803_),
    .B1(_06821_),
    .B2(_01178_),
    .ZN(_07001_));
 AOI221_X1 _24160_ (.A(_07001_),
    .B1(\alu_adder_result_ex[21] ),
    .B2(_03929_),
    .C1(\cs_registers_i.csr_mepc_o[21] ),
    .C2(_03923_),
    .ZN(_07002_));
 NAND2_X1 _24161_ (.A1(net23),
    .A2(_06889_),
    .ZN(_07003_));
 NAND2_X1 _24162_ (.A1(_07002_),
    .A2(_07003_),
    .ZN(_07004_));
 NAND2_X1 _24163_ (.A1(_03937_),
    .A2(_07004_),
    .ZN(_07005_));
 INV_X1 _24164_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .ZN(_07006_));
 OAI21_X2 _24165_ (.A(_07005_),
    .B1(_03937_),
    .B2(_07006_),
    .ZN(_07007_));
 NOR3_X2 _24166_ (.A1(_03957_),
    .A2(_06988_),
    .A3(_06995_),
    .ZN(_07008_));
 AOI21_X4 _24167_ (.A(_07008_),
    .B1(_04154_),
    .B2(_06981_),
    .ZN(_07009_));
 NAND3_X1 _24168_ (.A1(_06969_),
    .A2(_06984_),
    .A3(_07009_),
    .ZN(_07010_));
 XOR2_X1 _24169_ (.A(_07007_),
    .B(_07010_),
    .Z(_07011_));
 AOI21_X1 _24170_ (.A(_06999_),
    .B1(_07011_),
    .B2(_06880_),
    .ZN(_01353_));
 AOI22_X1 _24171_ (.A1(\cs_registers_i.csr_mepc_o[22] ),
    .A2(_03924_),
    .B1(_03927_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .ZN(_07012_));
 OAI21_X1 _24172_ (.A(_07012_),
    .B1(_06895_),
    .B2(_01179_),
    .ZN(_07013_));
 AOI21_X2 _24173_ (.A(_07013_),
    .B1(_06889_),
    .B2(net24),
    .ZN(_07014_));
 NAND2_X1 _24174_ (.A1(_03937_),
    .A2(_07014_),
    .ZN(_07015_));
 AOI21_X2 _24175_ (.A(_07015_),
    .B1(\alu_adder_result_ex[22] ),
    .B2(_03930_),
    .ZN(_07016_));
 NOR2_X1 _24176_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(_03937_),
    .ZN(_07017_));
 NOR2_X2 _24177_ (.A1(_07017_),
    .A2(_07016_),
    .ZN(_07018_));
 NAND4_X1 _24178_ (.A1(_06965_),
    .A2(_06983_),
    .A3(_07007_),
    .A4(_07009_),
    .ZN(_07019_));
 MUX2_X1 _24179_ (.A(_07016_),
    .B(_07018_),
    .S(_07019_),
    .Z(_07020_));
 NAND3_X1 _24180_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(_06858_),
    .A3(_04164_),
    .ZN(_07021_));
 NAND2_X1 _24181_ (.A1(_16107_),
    .A2(_07017_),
    .ZN(_07022_));
 OAI21_X1 _24182_ (.A(_07021_),
    .B1(_07022_),
    .B2(_07019_),
    .ZN(_07023_));
 OR2_X1 _24183_ (.A1(_07020_),
    .A2(_07023_),
    .ZN(_01354_));
 AOI22_X1 _24184_ (.A1(\cs_registers_i.csr_mepc_o[23] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .ZN(_07024_));
 OAI21_X1 _24185_ (.A(_07024_),
    .B1(_06895_),
    .B2(_01180_),
    .ZN(_07025_));
 AOI21_X2 _24186_ (.A(_07025_),
    .B1(_06889_),
    .B2(net25),
    .ZN(_07026_));
 NAND2_X1 _24187_ (.A1(_03937_),
    .A2(_07026_),
    .ZN(_07027_));
 AOI21_X1 _24188_ (.A(_07027_),
    .B1(\alu_adder_result_ex[23] ),
    .B2(_03930_),
    .ZN(_07028_));
 INV_X2 _24189_ (.A(_07028_),
    .ZN(_07029_));
 OAI21_X4 _24190_ (.A(_07029_),
    .B1(_03938_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .ZN(_07030_));
 NAND4_X1 _24191_ (.A1(_06984_),
    .A2(_07007_),
    .A3(_07009_),
    .A4(_07018_),
    .ZN(_07031_));
 NOR2_X1 _24192_ (.A1(_06930_),
    .A2(_07031_),
    .ZN(_07032_));
 XNOR2_X1 _24193_ (.A(_07030_),
    .B(_07032_),
    .ZN(_07033_));
 MUX2_X1 _24194_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .B(_07033_),
    .S(_06880_),
    .Z(_01355_));
 AOI22_X1 _24195_ (.A1(\cs_registers_i.csr_mepc_o[24] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .ZN(_07034_));
 OAI21_X1 _24196_ (.A(_07034_),
    .B1(_06895_),
    .B2(_01181_),
    .ZN(_07035_));
 AOI21_X2 _24197_ (.A(_07035_),
    .B1(_06889_),
    .B2(net26),
    .ZN(_07036_));
 NAND2_X1 _24198_ (.A1(_03936_),
    .A2(_07036_),
    .ZN(_07037_));
 AOI21_X2 _24199_ (.A(_07037_),
    .B1(\alu_adder_result_ex[24] ),
    .B2(_03930_),
    .ZN(_07038_));
 NOR2_X1 _24200_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(_03937_),
    .ZN(_07039_));
 OR2_X2 _24201_ (.A1(_07038_),
    .A2(_07039_),
    .ZN(_07040_));
 NAND2_X1 _24202_ (.A1(_06911_),
    .A2(_06929_),
    .ZN(_07041_));
 NOR3_X1 _24203_ (.A1(_07041_),
    .A2(_07030_),
    .A3(_07031_),
    .ZN(_07042_));
 XNOR2_X1 _24204_ (.A(_07040_),
    .B(_07042_),
    .ZN(_07043_));
 MUX2_X1 _24205_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .B(_07043_),
    .S(_06880_),
    .Z(_01356_));
 NAND3_X1 _24206_ (.A1(_03844_),
    .A2(_01182_),
    .A3(_06989_),
    .ZN(_07044_));
 OR3_X1 _24207_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_03878_),
    .A3(_03953_),
    .ZN(_07045_));
 NAND3_X1 _24208_ (.A1(_03893_),
    .A2(_07044_),
    .A3(_07045_),
    .ZN(_07046_));
 AOI22_X1 _24209_ (.A1(\cs_registers_i.csr_mepc_o[25] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .ZN(_07047_));
 NAND2_X1 _24210_ (.A1(_07046_),
    .A2(_07047_),
    .ZN(_07048_));
 AOI221_X2 _24211_ (.A(_07048_),
    .B1(\alu_adder_result_ex[25] ),
    .B2(_03930_),
    .C1(net27),
    .C2(_06888_),
    .ZN(_07049_));
 OR2_X4 _24212_ (.A1(_07049_),
    .A2(_04154_),
    .ZN(_07050_));
 INV_X1 _24213_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .ZN(_07051_));
 OAI21_X4 _24214_ (.A(_07050_),
    .B1(_03938_),
    .B2(_07051_),
    .ZN(_07052_));
 OR2_X1 _24215_ (.A1(_07017_),
    .A2(_07016_),
    .ZN(_07053_));
 NAND4_X2 _24216_ (.A1(_06964_),
    .A2(_06983_),
    .A3(_07007_),
    .A4(_07009_),
    .ZN(_07054_));
 NOR4_X4 _24217_ (.A1(_07053_),
    .A2(_07030_),
    .A3(_07054_),
    .A4(_07040_),
    .ZN(_07055_));
 NAND2_X2 _24218_ (.A1(_06969_),
    .A2(_07055_),
    .ZN(_07056_));
 XNOR2_X1 _24219_ (.A(_07052_),
    .B(_07056_),
    .ZN(_07057_));
 CLKBUF_X3 _24220_ (.A(_06879_),
    .Z(_07058_));
 MUX2_X1 _24221_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .B(_07057_),
    .S(_07058_),
    .Z(_01357_));
 NOR2_X2 _24222_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(_03938_),
    .ZN(_07059_));
 NAND2_X1 _24223_ (.A1(\cs_registers_i.csr_mepc_o[26] ),
    .A2(_03924_),
    .ZN(_07060_));
 OAI21_X1 _24224_ (.A(_07060_),
    .B1(_06895_),
    .B2(_01183_),
    .ZN(_07061_));
 AOI221_X2 _24225_ (.A(_07061_),
    .B1(_06888_),
    .B2(net28),
    .C1(\cs_registers_i.csr_depc_o[26] ),
    .C2(_03927_),
    .ZN(_07062_));
 AND2_X1 _24226_ (.A1(_03937_),
    .A2(_07062_),
    .ZN(_07063_));
 NAND2_X1 _24227_ (.A1(_03931_),
    .A2(\alu_adder_result_ex[26] ),
    .ZN(_07064_));
 AOI21_X4 _24228_ (.A(_07059_),
    .B1(_07063_),
    .B2(_07064_),
    .ZN(_07065_));
 AND3_X1 _24229_ (.A1(_06911_),
    .A2(_06929_),
    .A3(_07055_),
    .ZN(_07066_));
 NAND2_X1 _24230_ (.A1(_07052_),
    .A2(_07066_),
    .ZN(_07067_));
 XNOR2_X1 _24231_ (.A(_07065_),
    .B(_07067_),
    .ZN(_07068_));
 MUX2_X1 _24232_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .B(_07068_),
    .S(_07058_),
    .Z(_01358_));
 NAND3_X1 _24233_ (.A1(_03844_),
    .A2(_00007_),
    .A3(_06989_),
    .ZN(_07069_));
 OR3_X1 _24234_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_03878_),
    .A3(_03953_),
    .ZN(_07070_));
 NAND3_X1 _24235_ (.A1(_03893_),
    .A2(_07069_),
    .A3(_07070_),
    .ZN(_07071_));
 AOI22_X1 _24236_ (.A1(\cs_registers_i.csr_mepc_o[27] ),
    .A2(_03923_),
    .B1(_03926_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .ZN(_07072_));
 NAND2_X1 _24237_ (.A1(_07071_),
    .A2(_07072_),
    .ZN(_07073_));
 AOI221_X2 _24238_ (.A(_07073_),
    .B1(\alu_adder_result_ex[27] ),
    .B2(_03930_),
    .C1(net29),
    .C2(_06889_),
    .ZN(_07074_));
 OR2_X2 _24239_ (.A1(_07074_),
    .A2(_04154_),
    .ZN(_07075_));
 INV_X1 _24240_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .ZN(_07076_));
 OAI21_X2 _24241_ (.A(_07075_),
    .B1(_03938_),
    .B2(_07076_),
    .ZN(_07077_));
 NAND4_X1 _24242_ (.A1(_06969_),
    .A2(_07052_),
    .A3(_07055_),
    .A4(_07065_),
    .ZN(_07078_));
 XNOR2_X1 _24243_ (.A(_07077_),
    .B(_07078_),
    .ZN(_07079_));
 MUX2_X1 _24244_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .B(_07079_),
    .S(_07058_),
    .Z(_01359_));
 NAND3_X1 _24245_ (.A1(_03844_),
    .A2(_00008_),
    .A3(_06989_),
    .ZN(_07080_));
 OR3_X1 _24246_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_03878_),
    .A3(_06989_),
    .ZN(_07081_));
 NAND3_X1 _24247_ (.A1(_03893_),
    .A2(_07080_),
    .A3(_07081_),
    .ZN(_07082_));
 AOI22_X2 _24248_ (.A1(\cs_registers_i.csr_mepc_o[28] ),
    .A2(_03924_),
    .B1(_03927_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .ZN(_07083_));
 NAND2_X1 _24249_ (.A1(net30),
    .A2(_06889_),
    .ZN(_07084_));
 NAND4_X2 _24250_ (.A1(_03938_),
    .A2(_07082_),
    .A3(_07083_),
    .A4(_07084_),
    .ZN(_07085_));
 AOI21_X2 _24251_ (.A(_07085_),
    .B1(\alu_adder_result_ex[28] ),
    .B2(_03931_),
    .ZN(_07086_));
 NOR2_X1 _24252_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .A2(_03938_),
    .ZN(_07087_));
 NOR2_X1 _24253_ (.A1(_07086_),
    .A2(_07087_),
    .ZN(_07088_));
 NAND3_X1 _24254_ (.A1(_07052_),
    .A2(_07065_),
    .A3(_07077_),
    .ZN(_07089_));
 INV_X1 _24255_ (.A(_07089_),
    .ZN(_07090_));
 NAND2_X1 _24256_ (.A1(_07066_),
    .A2(_07090_),
    .ZN(_07091_));
 XNOR2_X1 _24257_ (.A(_07088_),
    .B(_07091_),
    .ZN(_07092_));
 MUX2_X1 _24258_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .B(_07092_),
    .S(_07058_),
    .Z(_01360_));
 AOI22_X2 _24259_ (.A1(\cs_registers_i.csr_mepc_o[29] ),
    .A2(_03924_),
    .B1(_03927_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .ZN(_07093_));
 OAI21_X2 _24260_ (.A(_07093_),
    .B1(_06895_),
    .B2(_00009_),
    .ZN(_07094_));
 AOI221_X2 _24261_ (.A(_07094_),
    .B1(\alu_adder_result_ex[29] ),
    .B2(_03930_),
    .C1(net31),
    .C2(_06889_),
    .ZN(_07095_));
 NOR2_X4 _24262_ (.A1(_07095_),
    .A2(_04154_),
    .ZN(_07096_));
 AOI21_X4 _24263_ (.A(_07096_),
    .B1(_06852_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .ZN(_07097_));
 OR2_X1 _24264_ (.A1(_07086_),
    .A2(_07087_),
    .ZN(_07098_));
 NOR3_X1 _24265_ (.A1(_07056_),
    .A2(_07098_),
    .A3(_07089_),
    .ZN(_07099_));
 XNOR2_X1 _24266_ (.A(_07097_),
    .B(_07099_),
    .ZN(_07100_));
 MUX2_X1 _24267_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .B(_07100_),
    .S(_07058_),
    .Z(_01361_));
 MUX2_X1 _24268_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .S(_07058_),
    .Z(_01362_));
 AOI22_X1 _24269_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_03924_),
    .B1(_03927_),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_07101_));
 OAI21_X1 _24270_ (.A(_07101_),
    .B1(_06895_),
    .B2(_00010_),
    .ZN(_07102_));
 AOI21_X2 _24271_ (.A(_07102_),
    .B1(_06889_),
    .B2(net32),
    .ZN(_07103_));
 NAND2_X1 _24272_ (.A1(_03938_),
    .A2(_07103_),
    .ZN(_07104_));
 AOI21_X4 _24273_ (.A(_07104_),
    .B1(\alu_adder_result_ex[30] ),
    .B2(_03931_),
    .ZN(_07105_));
 INV_X1 _24274_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .ZN(_07106_));
 AOI21_X2 _24275_ (.A(_07105_),
    .B1(_06852_),
    .B2(_07106_),
    .ZN(_07107_));
 NOR3_X1 _24276_ (.A1(_07098_),
    .A2(_07089_),
    .A3(_07097_),
    .ZN(_07108_));
 NAND2_X1 _24277_ (.A1(_07066_),
    .A2(_07108_),
    .ZN(_07109_));
 XNOR2_X1 _24278_ (.A(_07107_),
    .B(_07109_),
    .ZN(_07110_));
 MUX2_X1 _24279_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .B(_07110_),
    .S(_07058_),
    .Z(_01363_));
 NAND2_X1 _24280_ (.A1(_07107_),
    .A2(_07108_),
    .ZN(_07111_));
 NOR3_X1 _24281_ (.A1(_04164_),
    .A2(_07056_),
    .A3(_07111_),
    .ZN(_07112_));
 MUX2_X1 _24282_ (.A(_04164_),
    .B(_07112_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .Z(_07113_));
 NAND2_X1 _24283_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .A2(_06852_),
    .ZN(_07114_));
 NOR2_X1 _24284_ (.A1(_07056_),
    .A2(_07111_),
    .ZN(_07115_));
 AOI22_X2 _24285_ (.A1(\cs_registers_i.csr_mepc_o[31] ),
    .A2(_03924_),
    .B1(_03927_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .ZN(_07116_));
 OAI21_X2 _24286_ (.A(_07116_),
    .B1(_06895_),
    .B2(_00011_),
    .ZN(_07117_));
 AOI221_X2 _24287_ (.A(_07117_),
    .B1(_03931_),
    .B2(\alu_adder_result_ex[31] ),
    .C1(net33),
    .C2(_06889_),
    .ZN(_07118_));
 NOR2_X2 _24288_ (.A1(_07118_),
    .A2(_06852_),
    .ZN(_07119_));
 XNOR2_X1 _24289_ (.A(_07115_),
    .B(_07119_),
    .ZN(_07120_));
 AOI22_X1 _24290_ (.A1(_06863_),
    .A2(_07113_),
    .B1(_07114_),
    .B2(_07120_),
    .ZN(_01364_));
 MUX2_X1 _24291_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .S(_07058_),
    .Z(_01365_));
 XOR2_X1 _24292_ (.A(_16111_),
    .B(_06808_),
    .Z(_07121_));
 MUX2_X1 _24293_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .B(_07121_),
    .S(_07058_),
    .Z(_01366_));
 NAND3_X1 _24294_ (.A1(_16109_),
    .A2(_16110_),
    .A3(_06808_),
    .ZN(_07122_));
 XNOR2_X1 _24295_ (.A(_06818_),
    .B(_07122_),
    .ZN(_07123_));
 MUX2_X1 _24296_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .B(_07123_),
    .S(_07058_),
    .Z(_01367_));
 NOR2_X1 _24297_ (.A1(_06847_),
    .A2(_06848_),
    .ZN(_07124_));
 XNOR2_X1 _24298_ (.A(_07124_),
    .B(_06819_),
    .ZN(_07125_));
 MUX2_X1 _24299_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .B(_07125_),
    .S(_06879_),
    .Z(_01368_));
 NOR2_X1 _24300_ (.A1(_06840_),
    .A2(_06843_),
    .ZN(_07126_));
 NAND2_X1 _24301_ (.A1(_07124_),
    .A2(_06875_),
    .ZN(_07127_));
 XNOR2_X1 _24302_ (.A(_07126_),
    .B(_07127_),
    .ZN(_07128_));
 MUX2_X1 _24303_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .B(_07128_),
    .S(_06879_),
    .Z(_01369_));
 NAND4_X1 _24304_ (.A1(_16111_),
    .A2(_06808_),
    .A3(_06818_),
    .A4(_06849_),
    .ZN(_07129_));
 XNOR2_X1 _24305_ (.A(_06828_),
    .B(_07129_),
    .ZN(_07130_));
 MUX2_X1 _24306_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .B(_07130_),
    .S(_06879_),
    .Z(_01370_));
 NAND3_X1 _24307_ (.A1(_06828_),
    .A2(_06849_),
    .A3(_06875_),
    .ZN(_07131_));
 XNOR2_X1 _24308_ (.A(_06839_),
    .B(_07131_),
    .ZN(_07132_));
 MUX2_X1 _24309_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .B(_07132_),
    .S(_06879_),
    .Z(_01371_));
 BUF_X4 _24310_ (.A(_04158_),
    .Z(_07133_));
 BUF_X4 _24311_ (.A(_07133_),
    .Z(_07134_));
 MUX2_X1 _24312_ (.A(_03966_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .S(_07134_),
    .Z(_07135_));
 CLKBUF_X3 _24313_ (.A(_03979_),
    .Z(_07136_));
 BUF_X4 _24314_ (.A(_07136_),
    .Z(_07137_));
 INV_X2 _24315_ (.A(_04158_),
    .ZN(_07138_));
 NAND2_X1 _24316_ (.A1(_04155_),
    .A2(net134),
    .ZN(_07139_));
 NOR2_X1 _24317_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_07139_),
    .ZN(_07140_));
 NAND3_X2 _24318_ (.A1(_07137_),
    .A2(_07138_),
    .A3(_07140_),
    .ZN(_07141_));
 NAND2_X1 _24319_ (.A1(_00135_),
    .A2(_07141_),
    .ZN(_07142_));
 INV_X1 _24320_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .ZN(_07143_));
 INV_X1 _24321_ (.A(_07139_),
    .ZN(_07144_));
 NAND2_X2 _24322_ (.A1(_07143_),
    .A2(_07144_),
    .ZN(_07145_));
 NOR2_X1 _24323_ (.A1(_07137_),
    .A2(_07145_),
    .ZN(_07146_));
 NOR2_X1 _24324_ (.A1(_11422_),
    .A2(_06298_),
    .ZN(_07147_));
 AOI21_X1 _24325_ (.A(_11424_),
    .B1(_06303_),
    .B2(_06268_),
    .ZN(_07148_));
 OAI21_X2 _24326_ (.A(_07147_),
    .B1(_07148_),
    .B2(_11421_),
    .ZN(_07149_));
 AND2_X1 _24327_ (.A1(_00136_),
    .A2(_07145_),
    .ZN(_07150_));
 NAND2_X1 _24328_ (.A1(_03975_),
    .A2(_07150_),
    .ZN(_07151_));
 OAI21_X2 _24329_ (.A(_00135_),
    .B1(_07145_),
    .B2(_00136_),
    .ZN(_07152_));
 OAI21_X4 _24330_ (.A(_07151_),
    .B1(_07152_),
    .B2(_03975_),
    .ZN(_07153_));
 AOI21_X1 _24331_ (.A(_07153_),
    .B1(_03980_),
    .B2(_00137_),
    .ZN(_07154_));
 NAND3_X2 _24332_ (.A1(_06306_),
    .A2(_07149_),
    .A3(_07154_),
    .ZN(_07155_));
 OR2_X2 _24333_ (.A1(_06265_),
    .A2(_07155_),
    .ZN(_07156_));
 MUX2_X1 _24334_ (.A(_07142_),
    .B(_07146_),
    .S(_07156_),
    .Z(_07157_));
 BUF_X4 _24335_ (.A(_07157_),
    .Z(_07158_));
 BUF_X8 _24336_ (.A(_07158_),
    .Z(_07159_));
 MUX2_X1 _24337_ (.A(_03971_),
    .B(_07135_),
    .S(_07159_),
    .Z(_01372_));
 CLKBUF_X3 _24338_ (.A(_04156_),
    .Z(_07160_));
 MUX2_X1 _24339_ (.A(_03966_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(_07160_),
    .Z(_07161_));
 AOI21_X1 _24340_ (.A(_04156_),
    .B1(_07140_),
    .B2(_04158_),
    .ZN(_07162_));
 INV_X1 _24341_ (.A(_07162_),
    .ZN(_07163_));
 NOR3_X2 _24342_ (.A1(_06265_),
    .A2(_07155_),
    .A3(_07163_),
    .ZN(_07164_));
 AOI21_X4 _24343_ (.A(_07164_),
    .B1(_07141_),
    .B2(_07156_),
    .ZN(_07165_));
 CLKBUF_X3 _24344_ (.A(_07165_),
    .Z(_07166_));
 MUX2_X1 _24345_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B(_07161_),
    .S(_07166_),
    .Z(_01373_));
 NOR3_X4 _24346_ (.A1(_07138_),
    .A2(_04156_),
    .A3(_07145_),
    .ZN(_07167_));
 CLKBUF_X3 _24347_ (.A(_07167_),
    .Z(_07168_));
 MUX2_X1 _24348_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .B(_03966_),
    .S(_07168_),
    .Z(_01374_));
 INV_X2 _24349_ (.A(_03963_),
    .ZN(_07169_));
 BUF_X4 _24350_ (.A(_07169_),
    .Z(_07170_));
 NAND2_X1 _24351_ (.A1(_07170_),
    .A2(_06852_),
    .ZN(_07171_));
 NAND4_X4 _24352_ (.A1(_06253_),
    .A2(_06264_),
    .A3(_06306_),
    .A4(_07149_),
    .ZN(_07172_));
 NOR2_X1 _24353_ (.A1(_07150_),
    .A2(_07172_),
    .ZN(_07173_));
 AOI21_X1 _24354_ (.A(_07171_),
    .B1(_07173_),
    .B2(_03980_),
    .ZN(_07174_));
 NOR3_X1 _24355_ (.A1(_07170_),
    .A2(_03939_),
    .A3(_03974_),
    .ZN(_07175_));
 OAI22_X1 _24356_ (.A1(_16090_),
    .A2(_11426_),
    .B1(_06803_),
    .B2(_00554_),
    .ZN(_07176_));
 AOI21_X2 _24357_ (.A(_07176_),
    .B1(_06797_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .ZN(_07177_));
 AOI221_X1 _24358_ (.A(_07174_),
    .B1(_07175_),
    .B2(_07173_),
    .C1(_07177_),
    .C2(_06998_),
    .ZN(_01375_));
 BUF_X2 _24359_ (.A(\cs_registers_i.pc_if_i[11] ),
    .Z(_07178_));
 NOR2_X2 _24360_ (.A1(_07153_),
    .A2(_07172_),
    .ZN(_07179_));
 BUF_X4 _24361_ (.A(_07179_),
    .Z(_07180_));
 CLKBUF_X2 _24362_ (.A(\cs_registers_i.pc_if_i[3] ),
    .Z(_07181_));
 INV_X1 _24363_ (.A(_15355_),
    .ZN(_07182_));
 NAND2_X2 _24364_ (.A1(_07181_),
    .A2(_07182_),
    .ZN(_07183_));
 BUF_X2 _24365_ (.A(\cs_registers_i.pc_if_i[9] ),
    .Z(_07184_));
 CLKBUF_X2 _24366_ (.A(\cs_registers_i.pc_if_i[7] ),
    .Z(_07185_));
 CLKBUF_X2 _24367_ (.A(\cs_registers_i.pc_if_i[4] ),
    .Z(_07186_));
 CLKBUF_X2 _24368_ (.A(\cs_registers_i.pc_if_i[5] ),
    .Z(_07187_));
 AND3_X1 _24369_ (.A1(_07186_),
    .A2(_07187_),
    .A3(\cs_registers_i.pc_if_i[6] ),
    .ZN(_07188_));
 AND3_X1 _24370_ (.A1(_07185_),
    .A2(\cs_registers_i.pc_if_i[8] ),
    .A3(_07188_),
    .ZN(_07189_));
 NAND3_X2 _24371_ (.A1(_07184_),
    .A2(\cs_registers_i.pc_if_i[10] ),
    .A3(_07189_),
    .ZN(_07190_));
 NOR2_X1 _24372_ (.A1(_07183_),
    .A2(_07190_),
    .ZN(_07191_));
 AND4_X1 _24373_ (.A1(_07178_),
    .A2(_06905_),
    .A3(_07180_),
    .A4(_07191_),
    .ZN(_07192_));
 CLKBUF_X3 _24374_ (.A(_07179_),
    .Z(_07193_));
 NOR3_X1 _24375_ (.A1(_07178_),
    .A2(_06998_),
    .A3(_07193_),
    .ZN(_07194_));
 INV_X1 _24376_ (.A(_07178_),
    .ZN(_07195_));
 OAI21_X1 _24377_ (.A(_07195_),
    .B1(_07183_),
    .B2(_07190_),
    .ZN(_07196_));
 AOI21_X1 _24378_ (.A(_06870_),
    .B1(_07196_),
    .B2(_06858_),
    .ZN(_07197_));
 NOR3_X1 _24379_ (.A1(_07192_),
    .A2(_07194_),
    .A3(_07197_),
    .ZN(_01376_));
 NOR2_X1 _24380_ (.A1(_06858_),
    .A2(_06891_),
    .ZN(_07198_));
 CLKBUF_X2 _24381_ (.A(\cs_registers_i.pc_if_i[12] ),
    .Z(_07199_));
 CLKBUF_X3 _24382_ (.A(_07153_),
    .Z(_07200_));
 BUF_X4 _24383_ (.A(_07172_),
    .Z(_07201_));
 INV_X1 _24384_ (.A(_15833_),
    .ZN(_07202_));
 NOR2_X1 _24385_ (.A1(_07202_),
    .A2(_15354_),
    .ZN(_07203_));
 OAI21_X2 _24386_ (.A(_07181_),
    .B1(_15832_),
    .B2(_07203_),
    .ZN(_07204_));
 OR2_X1 _24387_ (.A1(_07190_),
    .A2(_07204_),
    .ZN(_07205_));
 NOR4_X1 _24388_ (.A1(_07195_),
    .A2(_07200_),
    .A3(_07201_),
    .A4(_07205_),
    .ZN(_07206_));
 XNOR2_X1 _24389_ (.A(_07199_),
    .B(_07206_),
    .ZN(_07207_));
 AOI21_X1 _24390_ (.A(_07198_),
    .B1(_07207_),
    .B2(_06863_),
    .ZN(_01377_));
 CLKBUF_X3 _24391_ (.A(_07153_),
    .Z(_07208_));
 CLKBUF_X3 _24392_ (.A(_07172_),
    .Z(_07209_));
 NAND3_X1 _24393_ (.A1(_07178_),
    .A2(_07199_),
    .A3(_07191_),
    .ZN(_07210_));
 NOR3_X1 _24394_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07210_),
    .ZN(_07211_));
 XNOR2_X1 _24395_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_07211_),
    .ZN(_07212_));
 AOI21_X1 _24396_ (.A(_06899_),
    .B1(_07212_),
    .B2(_06863_),
    .ZN(_01378_));
 INV_X1 _24397_ (.A(\cs_registers_i.pc_if_i[14] ),
    .ZN(_07213_));
 NAND3_X1 _24398_ (.A1(_07178_),
    .A2(_07199_),
    .A3(\cs_registers_i.pc_if_i[13] ),
    .ZN(_07214_));
 OR2_X1 _24399_ (.A1(_07205_),
    .A2(_07214_),
    .ZN(_07215_));
 CLKBUF_X3 _24400_ (.A(_07215_),
    .Z(_07216_));
 NAND2_X1 _24401_ (.A1(_06918_),
    .A2(_07216_),
    .ZN(_07217_));
 BUF_X4 _24402_ (.A(_07180_),
    .Z(_07218_));
 OAI21_X1 _24403_ (.A(_07217_),
    .B1(_07218_),
    .B2(_06998_),
    .ZN(_07219_));
 NOR4_X1 _24404_ (.A1(_07213_),
    .A2(_07200_),
    .A3(_07201_),
    .A4(_07216_),
    .ZN(_07220_));
 OR2_X1 _24405_ (.A1(_06998_),
    .A2(_07220_),
    .ZN(_07221_));
 AOI22_X1 _24406_ (.A1(_07213_),
    .A2(_07219_),
    .B1(_07221_),
    .B2(_06918_),
    .ZN(_01379_));
 BUF_X1 _24407_ (.A(\cs_registers_i.pc_if_i[15] ),
    .Z(_07222_));
 OR3_X2 _24408_ (.A1(_07183_),
    .A2(_07190_),
    .A3(_07214_),
    .ZN(_07223_));
 NOR4_X1 _24409_ (.A1(_07213_),
    .A2(_07153_),
    .A3(_07172_),
    .A4(_07223_),
    .ZN(_07224_));
 XNOR2_X1 _24410_ (.A(_07222_),
    .B(_07224_),
    .ZN(_07225_));
 OAI21_X1 _24411_ (.A(_06924_),
    .B1(_07225_),
    .B2(_06893_),
    .ZN(_01380_));
 NAND2_X1 _24412_ (.A1(\cs_registers_i.pc_if_i[14] ),
    .A2(_07222_),
    .ZN(_07226_));
 NOR4_X2 _24413_ (.A1(_07153_),
    .A2(_07172_),
    .A3(_07216_),
    .A4(_07226_),
    .ZN(_07227_));
 XNOR2_X1 _24414_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B(_07227_),
    .ZN(_07228_));
 BUF_X4 _24415_ (.A(_06858_),
    .Z(_07229_));
 AOI22_X1 _24416_ (.A1(_06939_),
    .A2(_06938_),
    .B1(_07228_),
    .B2(_07229_),
    .ZN(_01381_));
 INV_X1 _24417_ (.A(_06951_),
    .ZN(_07230_));
 INV_X1 _24418_ (.A(\cs_registers_i.pc_if_i[17] ),
    .ZN(_07231_));
 NAND3_X1 _24419_ (.A1(\cs_registers_i.pc_if_i[14] ),
    .A2(_07222_),
    .A3(\cs_registers_i.pc_if_i[16] ),
    .ZN(_07232_));
 NOR4_X1 _24420_ (.A1(_07153_),
    .A2(_07172_),
    .A3(_07223_),
    .A4(_07232_),
    .ZN(_07233_));
 XNOR2_X1 _24421_ (.A(_07231_),
    .B(_07233_),
    .ZN(_07234_));
 MUX2_X1 _24422_ (.A(_07230_),
    .B(_07234_),
    .S(_06858_),
    .Z(_01382_));
 CLKBUF_X2 _24423_ (.A(\cs_registers_i.pc_if_i[18] ),
    .Z(_07235_));
 NOR2_X1 _24424_ (.A1(_07231_),
    .A2(_07232_),
    .ZN(_07236_));
 INV_X1 _24425_ (.A(_07236_),
    .ZN(_07237_));
 NOR4_X1 _24426_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07216_),
    .A4(_07237_),
    .ZN(_07238_));
 XNOR2_X1 _24427_ (.A(_07235_),
    .B(_07238_),
    .ZN(_07239_));
 OAI21_X1 _24428_ (.A(_06959_),
    .B1(_07239_),
    .B2(_06893_),
    .ZN(_01383_));
 OR2_X2 _24429_ (.A1(_07153_),
    .A2(_07172_),
    .ZN(_07240_));
 BUF_X1 _24430_ (.A(\cs_registers_i.pc_if_i[19] ),
    .Z(_07241_));
 NAND3_X1 _24431_ (.A1(_07235_),
    .A2(_07241_),
    .A3(_07236_),
    .ZN(_07242_));
 NOR4_X1 _24432_ (.A1(_06975_),
    .A2(_07240_),
    .A3(_07223_),
    .A4(_07242_),
    .ZN(_07243_));
 NOR3_X1 _24433_ (.A1(_07241_),
    .A2(_06998_),
    .A3(_07180_),
    .ZN(_07244_));
 INV_X1 _24434_ (.A(_07241_),
    .ZN(_07245_));
 NAND2_X1 _24435_ (.A1(_07235_),
    .A2(_07236_),
    .ZN(_07246_));
 OAI21_X1 _24436_ (.A(_07245_),
    .B1(_07223_),
    .B2(_07246_),
    .ZN(_07247_));
 AOI21_X1 _24437_ (.A(_06975_),
    .B1(_07247_),
    .B2(_06858_),
    .ZN(_07248_));
 NOR3_X1 _24438_ (.A1(_07243_),
    .A2(_07244_),
    .A3(_07248_),
    .ZN(_01384_));
 CLKBUF_X2 _24439_ (.A(\cs_registers_i.pc_if_i[20] ),
    .Z(_07249_));
 NOR4_X2 _24440_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07216_),
    .A4(_07242_),
    .ZN(_07250_));
 XNOR2_X1 _24441_ (.A(_07249_),
    .B(_07250_),
    .ZN(_07251_));
 AOI21_X1 _24442_ (.A(_07008_),
    .B1(_07251_),
    .B2(_06863_),
    .ZN(_01385_));
 NOR3_X1 _24443_ (.A1(_15356_),
    .A2(_07208_),
    .A3(_07209_),
    .ZN(_07252_));
 BUF_X4 _24444_ (.A(_07240_),
    .Z(_07253_));
 AOI21_X1 _24445_ (.A(_07252_),
    .B1(_07253_),
    .B2(\cs_registers_i.pc_if_i[2] ),
    .ZN(_07254_));
 OAI21_X1 _24446_ (.A(_03934_),
    .B1(_07254_),
    .B2(_06893_),
    .ZN(_01386_));
 NOR2_X1 _24447_ (.A1(_07245_),
    .A2(_07246_),
    .ZN(_07255_));
 NAND2_X1 _24448_ (.A1(_07249_),
    .A2(_07255_),
    .ZN(_07256_));
 NOR4_X1 _24449_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07223_),
    .A4(_07256_),
    .ZN(_07257_));
 XNOR2_X1 _24450_ (.A(\cs_registers_i.pc_if_i[21] ),
    .B(_07257_),
    .ZN(_07258_));
 OAI21_X1 _24451_ (.A(_07005_),
    .B1(_07258_),
    .B2(_06893_),
    .ZN(_01387_));
 CLKBUF_X2 _24452_ (.A(\cs_registers_i.pc_if_i[22] ),
    .Z(_07259_));
 NAND3_X2 _24453_ (.A1(_07249_),
    .A2(\cs_registers_i.pc_if_i[21] ),
    .A3(_07255_),
    .ZN(_07260_));
 NOR4_X1 _24454_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07216_),
    .A4(_07260_),
    .ZN(_07261_));
 XNOR2_X1 _24455_ (.A(_07259_),
    .B(_07261_),
    .ZN(_07262_));
 AOI21_X1 _24456_ (.A(_07016_),
    .B1(_07262_),
    .B2(_06863_),
    .ZN(_01388_));
 BUF_X1 _24457_ (.A(\cs_registers_i.pc_if_i[23] ),
    .Z(_07263_));
 INV_X1 _24458_ (.A(_07259_),
    .ZN(_07264_));
 OR2_X1 _24459_ (.A1(_07223_),
    .A2(_07260_),
    .ZN(_07265_));
 NOR4_X1 _24460_ (.A1(_07264_),
    .A2(_07200_),
    .A3(_07201_),
    .A4(_07265_),
    .ZN(_07266_));
 XNOR2_X1 _24461_ (.A(_07263_),
    .B(_07266_),
    .ZN(_07267_));
 AOI21_X1 _24462_ (.A(_07028_),
    .B1(_07267_),
    .B2(_06863_),
    .ZN(_01389_));
 INV_X1 _24463_ (.A(_07260_),
    .ZN(_07268_));
 NAND3_X1 _24464_ (.A1(_07259_),
    .A2(_07263_),
    .A3(_07268_),
    .ZN(_07269_));
 NOR4_X1 _24465_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07216_),
    .A4(_07269_),
    .ZN(_07270_));
 XNOR2_X1 _24466_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B(_07270_),
    .ZN(_07271_));
 AOI21_X1 _24467_ (.A(_07038_),
    .B1(_07271_),
    .B2(_06863_),
    .ZN(_01390_));
 AND3_X1 _24468_ (.A1(_07259_),
    .A2(_07263_),
    .A3(\cs_registers_i.pc_if_i[24] ),
    .ZN(_07272_));
 NAND2_X1 _24469_ (.A1(\cs_registers_i.pc_if_i[25] ),
    .A2(_07272_),
    .ZN(_07273_));
 NOR2_X2 _24470_ (.A1(_07265_),
    .A2(_07273_),
    .ZN(_07274_));
 NAND3_X1 _24471_ (.A1(_07050_),
    .A2(_07193_),
    .A3(_07274_),
    .ZN(_07275_));
 OR3_X1 _24472_ (.A1(\cs_registers_i.pc_if_i[25] ),
    .A2(_03939_),
    .A3(_07179_),
    .ZN(_07276_));
 NOR2_X1 _24473_ (.A1(_07223_),
    .A2(_07260_),
    .ZN(_07277_));
 AOI21_X1 _24474_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B1(_07277_),
    .B2(_07272_),
    .ZN(_07278_));
 OAI21_X1 _24475_ (.A(_07050_),
    .B1(_07278_),
    .B2(_06998_),
    .ZN(_07279_));
 AND3_X1 _24476_ (.A1(_07275_),
    .A2(_07276_),
    .A3(_07279_),
    .ZN(_01391_));
 AND2_X1 _24477_ (.A1(_07064_),
    .A2(_07063_),
    .ZN(_07280_));
 CLKBUF_X2 _24478_ (.A(\cs_registers_i.pc_if_i[26] ),
    .Z(_07281_));
 OR3_X1 _24479_ (.A1(_07216_),
    .A2(_07260_),
    .A3(_07273_),
    .ZN(_07282_));
 NOR3_X1 _24480_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07282_),
    .ZN(_07283_));
 XNOR2_X1 _24481_ (.A(_07281_),
    .B(_07283_),
    .ZN(_07284_));
 AOI21_X1 _24482_ (.A(_07280_),
    .B1(_07284_),
    .B2(_06863_),
    .ZN(_01392_));
 BUF_X1 _24483_ (.A(\cs_registers_i.pc_if_i[27] ),
    .Z(_07285_));
 AND2_X1 _24484_ (.A1(_07281_),
    .A2(_07285_),
    .ZN(_07286_));
 NAND4_X1 _24485_ (.A1(_07075_),
    .A2(_07193_),
    .A3(_07274_),
    .A4(_07286_),
    .ZN(_07287_));
 OR3_X1 _24486_ (.A1(_07285_),
    .A2(_03939_),
    .A3(_07179_),
    .ZN(_07288_));
 AOI21_X1 _24487_ (.A(_07285_),
    .B1(_07274_),
    .B2(_07281_),
    .ZN(_07289_));
 OAI21_X1 _24488_ (.A(_07075_),
    .B1(_07289_),
    .B2(_06998_),
    .ZN(_07290_));
 AND3_X1 _24489_ (.A1(_07287_),
    .A2(_07288_),
    .A3(_07290_),
    .ZN(_01393_));
 NAND2_X1 _24490_ (.A1(_07281_),
    .A2(_07285_),
    .ZN(_07291_));
 NOR4_X1 _24491_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07282_),
    .A4(_07291_),
    .ZN(_07292_));
 XNOR2_X1 _24492_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(_07292_),
    .ZN(_07293_));
 AOI21_X1 _24493_ (.A(_07086_),
    .B1(_07293_),
    .B2(_07229_),
    .ZN(_01394_));
 INV_X1 _24494_ (.A(_07274_),
    .ZN(_07294_));
 AND2_X1 _24495_ (.A1(\cs_registers_i.pc_if_i[28] ),
    .A2(_07286_),
    .ZN(_07295_));
 NAND2_X1 _24496_ (.A1(\cs_registers_i.pc_if_i[29] ),
    .A2(_07295_),
    .ZN(_07296_));
 NOR4_X1 _24497_ (.A1(_07096_),
    .A2(_07253_),
    .A3(_07294_),
    .A4(_07296_),
    .ZN(_07297_));
 INV_X1 _24498_ (.A(_07096_),
    .ZN(_07298_));
 AOI21_X1 _24499_ (.A(\cs_registers_i.pc_if_i[29] ),
    .B1(_07274_),
    .B2(_07295_),
    .ZN(_07299_));
 OAI21_X1 _24500_ (.A(_07298_),
    .B1(_07299_),
    .B2(_06998_),
    .ZN(_07300_));
 OR2_X1 _24501_ (.A1(\cs_registers_i.pc_if_i[29] ),
    .A2(_03939_),
    .ZN(_07301_));
 OAI21_X1 _24502_ (.A(_07300_),
    .B1(_07301_),
    .B2(_07218_),
    .ZN(_07302_));
 NOR2_X1 _24503_ (.A1(_07297_),
    .A2(_07302_),
    .ZN(_01395_));
 NOR4_X1 _24504_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07282_),
    .A4(_07296_),
    .ZN(_07303_));
 XNOR2_X1 _24505_ (.A(\cs_registers_i.pc_if_i[30] ),
    .B(_07303_),
    .ZN(_07304_));
 AOI21_X1 _24506_ (.A(_07105_),
    .B1(_07304_),
    .B2(_07229_),
    .ZN(_01396_));
 NOR3_X1 _24507_ (.A1(_15355_),
    .A2(_07208_),
    .A3(_07209_),
    .ZN(_07305_));
 XNOR2_X1 _24508_ (.A(_07181_),
    .B(_07305_),
    .ZN(_07306_));
 AOI21_X1 _24509_ (.A(_03956_),
    .B1(_07306_),
    .B2(_07229_),
    .ZN(_01397_));
 INV_X2 _24510_ (.A(_07119_),
    .ZN(_07307_));
 INV_X1 _24511_ (.A(\cs_registers_i.pc_if_i[30] ),
    .ZN(_07308_));
 NOR3_X1 _24512_ (.A1(_07308_),
    .A2(_07294_),
    .A3(_07296_),
    .ZN(_07309_));
 NAND2_X1 _24513_ (.A1(\cs_registers_i.pc_if_i[31] ),
    .A2(_07309_),
    .ZN(_07310_));
 OAI21_X1 _24514_ (.A(_06858_),
    .B1(_07253_),
    .B2(_07310_),
    .ZN(_07311_));
 OAI22_X1 _24515_ (.A1(_06998_),
    .A2(_07193_),
    .B1(_07309_),
    .B2(_07119_),
    .ZN(_07312_));
 INV_X1 _24516_ (.A(\cs_registers_i.pc_if_i[31] ),
    .ZN(_07313_));
 AOI22_X1 _24517_ (.A1(_07307_),
    .A2(_07311_),
    .B1(_07312_),
    .B2(_07313_),
    .ZN(_01398_));
 NOR3_X1 _24518_ (.A1(_07208_),
    .A2(_07209_),
    .A3(_07204_),
    .ZN(_07314_));
 XNOR2_X1 _24519_ (.A(_07186_),
    .B(_07314_),
    .ZN(_07315_));
 AOI21_X1 _24520_ (.A(_06806_),
    .B1(_07315_),
    .B2(_07229_),
    .ZN(_01399_));
 INV_X1 _24521_ (.A(_07186_),
    .ZN(_07316_));
 NOR4_X2 _24522_ (.A1(_07316_),
    .A2(_07153_),
    .A3(_07172_),
    .A4(_07183_),
    .ZN(_07317_));
 XNOR2_X1 _24523_ (.A(_07187_),
    .B(_07317_),
    .ZN(_07318_));
 AOI21_X1 _24524_ (.A(_06816_),
    .B1(_07318_),
    .B2(_07229_),
    .ZN(_01400_));
 NAND2_X1 _24525_ (.A1(_07186_),
    .A2(_07187_),
    .ZN(_07319_));
 NOR4_X1 _24526_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07319_),
    .A4(_07204_),
    .ZN(_07320_));
 XNOR2_X1 _24527_ (.A(\cs_registers_i.pc_if_i[6] ),
    .B(_07320_),
    .ZN(_07321_));
 AOI21_X1 _24528_ (.A(_06847_),
    .B1(_07321_),
    .B2(_07229_),
    .ZN(_01401_));
 INV_X1 _24529_ (.A(_07188_),
    .ZN(_07322_));
 NOR4_X1 _24530_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07183_),
    .A4(_07322_),
    .ZN(_07323_));
 XNOR2_X1 _24531_ (.A(_07185_),
    .B(_07323_),
    .ZN(_07324_));
 AOI21_X1 _24532_ (.A(_06843_),
    .B1(_07324_),
    .B2(_07229_),
    .ZN(_01402_));
 NAND2_X1 _24533_ (.A1(_07185_),
    .A2(_07188_),
    .ZN(_07325_));
 NOR4_X1 _24534_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07325_),
    .A4(_07204_),
    .ZN(_07326_));
 XNOR2_X1 _24535_ (.A(\cs_registers_i.pc_if_i[8] ),
    .B(_07326_),
    .ZN(_07327_));
 AOI21_X1 _24536_ (.A(_06826_),
    .B1(_07327_),
    .B2(_07229_),
    .ZN(_01403_));
 INV_X1 _24537_ (.A(_07189_),
    .ZN(_07328_));
 NOR4_X1 _24538_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07183_),
    .A4(_07328_),
    .ZN(_07329_));
 XNOR2_X1 _24539_ (.A(_07184_),
    .B(_07329_),
    .ZN(_07330_));
 OAI21_X1 _24540_ (.A(_06837_),
    .B1(_07330_),
    .B2(_06893_),
    .ZN(_01404_));
 NAND2_X1 _24541_ (.A1(_07184_),
    .A2(_07189_),
    .ZN(_07331_));
 NOR4_X1 _24542_ (.A1(_07200_),
    .A2(_07201_),
    .A3(_07331_),
    .A4(_07204_),
    .ZN(_07332_));
 XNOR2_X1 _24543_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(_07332_),
    .ZN(_07333_));
 OAI21_X1 _24544_ (.A(_06856_),
    .B1(_07333_),
    .B2(_06893_),
    .ZN(_01405_));
 MUX2_X1 _24545_ (.A(net104),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_07334_));
 MUX2_X1 _24546_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B(_07334_),
    .S(_07159_),
    .Z(_01406_));
 MUX2_X1 _24547_ (.A(net105),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(_04157_),
    .Z(_07335_));
 MUX2_X1 _24548_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .B(_07335_),
    .S(_07159_),
    .Z(_01407_));
 MUX2_X1 _24549_ (.A(net106),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(_04157_),
    .Z(_07336_));
 MUX2_X1 _24550_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .B(_07336_),
    .S(_07159_),
    .Z(_01408_));
 MUX2_X1 _24551_ (.A(net107),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(_04157_),
    .Z(_07337_));
 MUX2_X1 _24552_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .B(_07337_),
    .S(_07159_),
    .Z(_01409_));
 MUX2_X1 _24553_ (.A(net108),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(_04157_),
    .Z(_07338_));
 MUX2_X1 _24554_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .B(_07338_),
    .S(_07159_),
    .Z(_01410_));
 MUX2_X1 _24555_ (.A(net109),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(_04157_),
    .Z(_07339_));
 MUX2_X1 _24556_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .B(_07339_),
    .S(_07159_),
    .Z(_01411_));
 MUX2_X1 _24557_ (.A(net110),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(_04158_),
    .Z(_07340_));
 MUX2_X1 _24558_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .B(_07340_),
    .S(_07159_),
    .Z(_01412_));
 MUX2_X1 _24559_ (.A(_03968_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(_07134_),
    .Z(_07341_));
 MUX2_X1 _24560_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .B(_07341_),
    .S(_07159_),
    .Z(_01413_));
 MUX2_X1 _24561_ (.A(_03967_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(_07134_),
    .Z(_07342_));
 MUX2_X1 _24562_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .B(_07342_),
    .S(_07159_),
    .Z(_01414_));
 MUX2_X1 _24563_ (.A(net111),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(_07134_),
    .Z(_07343_));
 BUF_X8 _24564_ (.A(_07158_),
    .Z(_07344_));
 MUX2_X1 _24565_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .B(_07343_),
    .S(_07344_),
    .Z(_01415_));
 MUX2_X1 _24566_ (.A(net112),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(_07134_),
    .Z(_07345_));
 MUX2_X1 _24567_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .B(_07345_),
    .S(_07344_),
    .Z(_01416_));
 MUX2_X1 _24568_ (.A(net113),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(_04157_),
    .Z(_07346_));
 MUX2_X1 _24569_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B(_07346_),
    .S(_07344_),
    .Z(_01417_));
 MUX2_X1 _24570_ (.A(net114),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(_07134_),
    .Z(_07347_));
 MUX2_X1 _24571_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .B(_07347_),
    .S(_07344_),
    .Z(_01418_));
 MUX2_X1 _24572_ (.A(net115),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(_07134_),
    .Z(_07348_));
 MUX2_X1 _24573_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .B(_07348_),
    .S(_07344_),
    .Z(_01419_));
 MUX2_X1 _24574_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(_07134_),
    .Z(_07349_));
 MUX2_X1 _24575_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .B(_07349_),
    .S(_07344_),
    .Z(_01420_));
 MUX2_X1 _24576_ (.A(net117),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(_07134_),
    .Z(_07350_));
 MUX2_X1 _24577_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .B(_07350_),
    .S(_07344_),
    .Z(_01421_));
 MUX2_X1 _24578_ (.A(net118),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(_07134_),
    .Z(_07351_));
 MUX2_X1 _24579_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .B(_07351_),
    .S(_07344_),
    .Z(_01422_));
 MUX2_X1 _24580_ (.A(net119),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(_07133_),
    .Z(_07352_));
 MUX2_X1 _24581_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .B(_07352_),
    .S(_07344_),
    .Z(_01423_));
 MUX2_X1 _24582_ (.A(net120),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(_07133_),
    .Z(_07353_));
 MUX2_X1 _24583_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .B(_07353_),
    .S(_07344_),
    .Z(_01424_));
 MUX2_X1 _24584_ (.A(net121),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(_07133_),
    .Z(_07354_));
 BUF_X8 _24585_ (.A(_07158_),
    .Z(_07355_));
 MUX2_X1 _24586_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .B(_07354_),
    .S(_07355_),
    .Z(_01425_));
 MUX2_X1 _24587_ (.A(net122),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(_07133_),
    .Z(_07356_));
 MUX2_X1 _24588_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .B(_07356_),
    .S(_07355_),
    .Z(_01426_));
 MUX2_X1 _24589_ (.A(net123),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(_07133_),
    .Z(_07357_));
 MUX2_X1 _24590_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .B(_07357_),
    .S(_07355_),
    .Z(_01427_));
 MUX2_X1 _24591_ (.A(net124),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(_04157_),
    .Z(_07358_));
 MUX2_X1 _24592_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .B(_07358_),
    .S(_07355_),
    .Z(_01428_));
 MUX2_X1 _24593_ (.A(net125),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(_07133_),
    .Z(_07359_));
 MUX2_X1 _24594_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .B(_07359_),
    .S(_07355_),
    .Z(_01429_));
 MUX2_X1 _24595_ (.A(net126),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(_07133_),
    .Z(_07360_));
 MUX2_X1 _24596_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .B(_07360_),
    .S(_07355_),
    .Z(_01430_));
 MUX2_X1 _24597_ (.A(net104),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(_07160_),
    .Z(_07361_));
 MUX2_X1 _24598_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .B(_07361_),
    .S(_07166_),
    .Z(_01431_));
 MUX2_X1 _24599_ (.A(net113),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(_07160_),
    .Z(_07362_));
 MUX2_X1 _24600_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .B(_07362_),
    .S(_07166_),
    .Z(_01432_));
 MUX2_X1 _24601_ (.A(net124),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(_07160_),
    .Z(_07363_));
 MUX2_X1 _24602_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .B(_07363_),
    .S(_07166_),
    .Z(_01433_));
 MUX2_X1 _24603_ (.A(net127),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(_07160_),
    .Z(_07364_));
 MUX2_X1 _24604_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .B(_07364_),
    .S(_07166_),
    .Z(_01434_));
 MUX2_X1 _24605_ (.A(net128),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(_07160_),
    .Z(_07365_));
 MUX2_X1 _24606_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .B(_07365_),
    .S(_07166_),
    .Z(_01435_));
 MUX2_X1 _24607_ (.A(net129),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(_07160_),
    .Z(_07366_));
 MUX2_X1 _24608_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .B(_07366_),
    .S(_07166_),
    .Z(_01436_));
 MUX2_X1 _24609_ (.A(net130),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(_07160_),
    .Z(_07367_));
 MUX2_X1 _24610_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .B(_07367_),
    .S(_07166_),
    .Z(_01437_));
 MUX2_X1 _24611_ (.A(net131),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(_07160_),
    .Z(_07368_));
 MUX2_X1 _24612_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .B(_07368_),
    .S(_07166_),
    .Z(_01438_));
 MUX2_X1 _24613_ (.A(net127),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(_04158_),
    .Z(_07369_));
 MUX2_X1 _24614_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .B(_07369_),
    .S(_07355_),
    .Z(_01439_));
 MUX2_X1 _24615_ (.A(net132),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(_07160_),
    .Z(_07370_));
 MUX2_X1 _24616_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .B(_07370_),
    .S(_07166_),
    .Z(_01440_));
 CLKBUF_X3 _24617_ (.A(_04156_),
    .Z(_07371_));
 MUX2_X1 _24618_ (.A(net133),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(_07371_),
    .Z(_07372_));
 CLKBUF_X3 _24619_ (.A(_07165_),
    .Z(_07373_));
 MUX2_X1 _24620_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .B(_07372_),
    .S(_07373_),
    .Z(_01441_));
 MUX2_X1 _24621_ (.A(net105),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(_07371_),
    .Z(_07374_));
 MUX2_X1 _24622_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .B(_07374_),
    .S(_07373_),
    .Z(_01442_));
 MUX2_X1 _24623_ (.A(net106),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(_07371_),
    .Z(_07375_));
 MUX2_X1 _24624_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .B(_07375_),
    .S(_07373_),
    .Z(_01443_));
 MUX2_X1 _24625_ (.A(net107),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(_07371_),
    .Z(_07376_));
 MUX2_X1 _24626_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .B(_07376_),
    .S(_07373_),
    .Z(_01444_));
 MUX2_X1 _24627_ (.A(net108),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(_07371_),
    .Z(_07377_));
 MUX2_X1 _24628_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .B(_07377_),
    .S(_07373_),
    .Z(_01445_));
 MUX2_X1 _24629_ (.A(net109),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(_07371_),
    .Z(_07378_));
 MUX2_X1 _24630_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .B(_07378_),
    .S(_07373_),
    .Z(_01446_));
 MUX2_X1 _24631_ (.A(net110),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(_07371_),
    .Z(_07379_));
 MUX2_X1 _24632_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .B(_07379_),
    .S(_07373_),
    .Z(_01447_));
 MUX2_X1 _24633_ (.A(_03968_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(_07371_),
    .Z(_07380_));
 MUX2_X1 _24634_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .B(_07380_),
    .S(_07373_),
    .Z(_01448_));
 MUX2_X1 _24635_ (.A(_03967_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(_07371_),
    .Z(_07381_));
 MUX2_X1 _24636_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .B(_07381_),
    .S(_07373_),
    .Z(_01449_));
 MUX2_X1 _24637_ (.A(net128),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(_04157_),
    .Z(_07382_));
 MUX2_X1 _24638_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .B(_07382_),
    .S(_07355_),
    .Z(_01450_));
 MUX2_X1 _24639_ (.A(net111),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(_07371_),
    .Z(_07383_));
 MUX2_X1 _24640_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .B(_07383_),
    .S(_07373_),
    .Z(_01451_));
 CLKBUF_X3 _24641_ (.A(_04156_),
    .Z(_07384_));
 MUX2_X1 _24642_ (.A(net112),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(_07384_),
    .Z(_07385_));
 CLKBUF_X3 _24643_ (.A(_07165_),
    .Z(_07386_));
 MUX2_X1 _24644_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .B(_07385_),
    .S(_07386_),
    .Z(_01452_));
 MUX2_X1 _24645_ (.A(net114),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(_07384_),
    .Z(_07387_));
 MUX2_X1 _24646_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .B(_07387_),
    .S(_07386_),
    .Z(_01453_));
 MUX2_X1 _24647_ (.A(net115),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(_07384_),
    .Z(_07388_));
 MUX2_X1 _24648_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .B(_07388_),
    .S(_07386_),
    .Z(_01454_));
 MUX2_X1 _24649_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(_07384_),
    .Z(_07389_));
 MUX2_X1 _24650_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .B(_07389_),
    .S(_07386_),
    .Z(_01455_));
 MUX2_X1 _24651_ (.A(net117),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(_07384_),
    .Z(_07390_));
 MUX2_X1 _24652_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .B(_07390_),
    .S(_07386_),
    .Z(_01456_));
 MUX2_X1 _24653_ (.A(net118),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(_07384_),
    .Z(_07391_));
 MUX2_X1 _24654_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .B(_07391_),
    .S(_07386_),
    .Z(_01457_));
 MUX2_X1 _24655_ (.A(net119),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(_07384_),
    .Z(_07392_));
 MUX2_X1 _24656_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .B(_07392_),
    .S(_07386_),
    .Z(_01458_));
 MUX2_X1 _24657_ (.A(net120),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(_07384_),
    .Z(_07393_));
 MUX2_X1 _24658_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .B(_07393_),
    .S(_07386_),
    .Z(_01459_));
 MUX2_X1 _24659_ (.A(net121),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(_07384_),
    .Z(_07394_));
 MUX2_X1 _24660_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .B(_07394_),
    .S(_07386_),
    .Z(_01460_));
 MUX2_X1 _24661_ (.A(net129),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(_04158_),
    .Z(_07395_));
 MUX2_X1 _24662_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .B(_07395_),
    .S(_07355_),
    .Z(_01461_));
 MUX2_X1 _24663_ (.A(net122),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(_07384_),
    .Z(_07396_));
 MUX2_X1 _24664_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .B(_07396_),
    .S(_07386_),
    .Z(_01462_));
 MUX2_X1 _24665_ (.A(net123),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(_04156_),
    .Z(_07397_));
 MUX2_X1 _24666_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .B(_07397_),
    .S(_07165_),
    .Z(_01463_));
 MUX2_X1 _24667_ (.A(net125),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(_04156_),
    .Z(_07398_));
 MUX2_X1 _24668_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .B(_07398_),
    .S(_07165_),
    .Z(_01464_));
 MUX2_X1 _24669_ (.A(net126),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(_04156_),
    .Z(_07399_));
 MUX2_X1 _24670_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .B(_07399_),
    .S(_07165_),
    .Z(_01465_));
 MUX2_X1 _24671_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .B(net104),
    .S(_07168_),
    .Z(_01466_));
 MUX2_X1 _24672_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .B(net113),
    .S(_07168_),
    .Z(_01467_));
 MUX2_X1 _24673_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .B(net124),
    .S(_07168_),
    .Z(_01468_));
 MUX2_X1 _24674_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .B(net127),
    .S(_07168_),
    .Z(_01469_));
 MUX2_X1 _24675_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .B(net128),
    .S(_07168_),
    .Z(_01470_));
 MUX2_X1 _24676_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .B(net129),
    .S(_07168_),
    .Z(_01471_));
 MUX2_X1 _24677_ (.A(net130),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_07400_));
 MUX2_X1 _24678_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .B(_07400_),
    .S(_07355_),
    .Z(_01472_));
 MUX2_X1 _24679_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .B(net130),
    .S(_07168_),
    .Z(_01473_));
 MUX2_X1 _24680_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .B(net131),
    .S(_07168_),
    .Z(_01474_));
 MUX2_X1 _24681_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .B(net132),
    .S(_07168_),
    .Z(_01475_));
 CLKBUF_X3 _24682_ (.A(_07167_),
    .Z(_07401_));
 MUX2_X1 _24683_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .B(net133),
    .S(_07401_),
    .Z(_01476_));
 MUX2_X1 _24684_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .B(net105),
    .S(_07401_),
    .Z(_01477_));
 MUX2_X1 _24685_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .B(net106),
    .S(_07401_),
    .Z(_01478_));
 MUX2_X1 _24686_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .B(net107),
    .S(_07401_),
    .Z(_01479_));
 MUX2_X1 _24687_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .B(net108),
    .S(_07401_),
    .Z(_01480_));
 MUX2_X1 _24688_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .B(net109),
    .S(_07401_),
    .Z(_01481_));
 MUX2_X1 _24689_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .B(net110),
    .S(_07401_),
    .Z(_01482_));
 MUX2_X1 _24690_ (.A(net131),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(_04158_),
    .Z(_07402_));
 MUX2_X1 _24691_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .B(_07402_),
    .S(_07158_),
    .Z(_01483_));
 MUX2_X1 _24692_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .B(_03968_),
    .S(_07401_),
    .Z(_01484_));
 MUX2_X1 _24693_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .B(_03967_),
    .S(_07401_),
    .Z(_01485_));
 MUX2_X1 _24694_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .B(net111),
    .S(_07401_),
    .Z(_01486_));
 CLKBUF_X3 _24695_ (.A(_07167_),
    .Z(_07403_));
 MUX2_X1 _24696_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .B(net112),
    .S(_07403_),
    .Z(_01487_));
 MUX2_X1 _24697_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .B(net114),
    .S(_07403_),
    .Z(_01488_));
 MUX2_X1 _24698_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .B(net115),
    .S(_07403_),
    .Z(_01489_));
 MUX2_X1 _24699_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .B(net116),
    .S(_07403_),
    .Z(_01490_));
 MUX2_X1 _24700_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .B(net117),
    .S(_07403_),
    .Z(_01491_));
 MUX2_X1 _24701_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .B(net118),
    .S(_07403_),
    .Z(_01492_));
 MUX2_X1 _24702_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .B(net119),
    .S(_07403_),
    .Z(_01493_));
 MUX2_X1 _24703_ (.A(net132),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(_04157_),
    .Z(_07404_));
 MUX2_X1 _24704_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .B(_07404_),
    .S(_07158_),
    .Z(_01494_));
 MUX2_X1 _24705_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .B(net120),
    .S(_07403_),
    .Z(_01495_));
 MUX2_X1 _24706_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .B(net121),
    .S(_07403_),
    .Z(_01496_));
 MUX2_X1 _24707_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .B(net122),
    .S(_07403_),
    .Z(_01497_));
 MUX2_X1 _24708_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .B(net123),
    .S(_07167_),
    .Z(_01498_));
 MUX2_X1 _24709_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .B(net125),
    .S(_07167_),
    .Z(_01499_));
 MUX2_X1 _24710_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .B(net126),
    .S(_07167_),
    .Z(_01500_));
 MUX2_X1 _24711_ (.A(net133),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(_04158_),
    .Z(_07405_));
 MUX2_X1 _24712_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .B(_07405_),
    .S(_07158_),
    .Z(_01501_));
 INV_X1 _24713_ (.A(_03959_),
    .ZN(_07406_));
 CLKBUF_X3 _24714_ (.A(_07406_),
    .Z(_07407_));
 NOR2_X1 _24715_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .A2(_07407_),
    .ZN(_07408_));
 AOI21_X1 _24716_ (.A(_07408_),
    .B1(_06872_),
    .B2(_07407_),
    .ZN(net224));
 NOR2_X1 _24717_ (.A1(net103),
    .A2(_04164_),
    .ZN(_07409_));
 CLKBUF_X3 _24718_ (.A(_07409_),
    .Z(_07410_));
 MUX2_X1 _24719_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .B(net224),
    .S(_07410_),
    .Z(_01502_));
 MUX2_X1 _24720_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .B(_06907_),
    .S(_07407_),
    .Z(net225));
 MUX2_X1 _24721_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .B(net225),
    .S(_07410_),
    .Z(_01503_));
 NAND2_X1 _24722_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .A2(_03959_),
    .ZN(_07411_));
 OAI21_X1 _24723_ (.A(_07411_),
    .B1(_06904_),
    .B2(_03959_),
    .ZN(net226));
 MUX2_X1 _24724_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .B(net226),
    .S(_07410_),
    .Z(_01504_));
 MUX2_X1 _24725_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .B(_06928_),
    .S(_07407_),
    .Z(net227));
 MUX2_X1 _24726_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .B(net227),
    .S(_07410_),
    .Z(_01505_));
 MUX2_X1 _24727_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .B(_06929_),
    .S(_07407_),
    .Z(net228));
 MUX2_X1 _24728_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .B(net228),
    .S(_07410_),
    .Z(_01506_));
 MUX2_X1 _24729_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .B(_06926_),
    .S(_07407_),
    .Z(net229));
 MUX2_X1 _24730_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .B(net229),
    .S(_07410_),
    .Z(_01507_));
 CLKBUF_X3 _24731_ (.A(_07406_),
    .Z(_07412_));
 MUX2_X1 _24732_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .B(_06940_),
    .S(_07412_),
    .Z(net230));
 MUX2_X1 _24733_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .B(net230),
    .S(_07410_),
    .Z(_01508_));
 MUX2_X1 _24734_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .B(_06963_),
    .S(_07412_),
    .Z(net231));
 MUX2_X1 _24735_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .B(net231),
    .S(_07410_),
    .Z(_01509_));
 MUX2_X1 _24736_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .B(_06961_),
    .S(_07412_),
    .Z(net232));
 MUX2_X1 _24737_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .B(net232),
    .S(_07410_),
    .Z(_01510_));
 OAI21_X1 _24738_ (.A(_07407_),
    .B1(_06967_),
    .B2(_06975_),
    .ZN(_07413_));
 INV_X1 _24739_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .ZN(_07414_));
 OAI21_X1 _24740_ (.A(_07413_),
    .B1(_07407_),
    .B2(_07414_),
    .ZN(net233));
 MUX2_X1 _24741_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .B(net233),
    .S(_07410_),
    .Z(_01511_));
 MUX2_X1 _24742_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .B(_07009_),
    .S(_07412_),
    .Z(net234));
 CLKBUF_X3 _24743_ (.A(_07409_),
    .Z(_07415_));
 MUX2_X1 _24744_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .B(net234),
    .S(_07415_),
    .Z(_01512_));
 MUX2_X1 _24745_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .B(_07007_),
    .S(_07412_),
    .Z(net235));
 MUX2_X1 _24746_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .B(net235),
    .S(_07415_),
    .Z(_01513_));
 MUX2_X1 _24747_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .B(_07018_),
    .S(_07412_),
    .Z(net236));
 MUX2_X1 _24748_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .B(net236),
    .S(_07415_),
    .Z(_01514_));
 NAND2_X1 _24749_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .A2(_03959_),
    .ZN(_07416_));
 OAI21_X2 _24750_ (.A(_07416_),
    .B1(_07030_),
    .B2(_03959_),
    .ZN(net237));
 MUX2_X1 _24751_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .B(net237),
    .S(_07415_),
    .Z(_01515_));
 NAND2_X1 _24752_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .A2(_03959_),
    .ZN(_07417_));
 OAI21_X1 _24753_ (.A(_07417_),
    .B1(_07040_),
    .B2(_03959_),
    .ZN(net238));
 MUX2_X1 _24754_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .B(net238),
    .S(_07415_),
    .Z(_01516_));
 MUX2_X1 _24755_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .B(_07052_),
    .S(_07412_),
    .Z(net239));
 MUX2_X1 _24756_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .B(net239),
    .S(_07415_),
    .Z(_01517_));
 MUX2_X1 _24757_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .B(_07065_),
    .S(_07412_),
    .Z(net240));
 MUX2_X1 _24758_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .B(net240),
    .S(_07415_),
    .Z(_01518_));
 MUX2_X1 _24759_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .B(_07077_),
    .S(_07412_),
    .Z(net241));
 MUX2_X1 _24760_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .B(net241),
    .S(_07415_),
    .Z(_01519_));
 MUX2_X1 _24761_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .B(_07088_),
    .S(_07412_),
    .Z(net242));
 MUX2_X1 _24762_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .B(net242),
    .S(_07415_),
    .Z(_01520_));
 NOR2_X1 _24763_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .A2(_07407_),
    .ZN(_07418_));
 AOI21_X2 _24764_ (.A(_07418_),
    .B1(_07097_),
    .B2(_07407_),
    .ZN(net243));
 MUX2_X1 _24765_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .B(net243),
    .S(_07415_),
    .Z(_01521_));
 CLKBUF_X3 _24766_ (.A(_07406_),
    .Z(_07419_));
 MUX2_X1 _24767_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .B(_16108_),
    .S(_07419_),
    .Z(net244));
 CLKBUF_X3 _24768_ (.A(_07409_),
    .Z(_07420_));
 MUX2_X1 _24769_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .B(net244),
    .S(_07420_),
    .Z(_01522_));
 MUX2_X1 _24770_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .B(_07107_),
    .S(_07419_),
    .Z(net245));
 MUX2_X1 _24771_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .B(net245),
    .S(_07420_),
    .Z(_01523_));
 NAND2_X2 _24772_ (.A1(_07307_),
    .A2(_07114_),
    .ZN(_07421_));
 MUX2_X1 _24773_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .B(_07421_),
    .S(_07419_),
    .Z(net246));
 MUX2_X1 _24774_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .B(net246),
    .S(_07420_),
    .Z(_01524_));
 MUX2_X1 _24775_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .B(_16110_),
    .S(_07419_),
    .Z(net247));
 MUX2_X1 _24776_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .B(net247),
    .S(_07420_),
    .Z(_01525_));
 MUX2_X1 _24777_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .B(_06808_),
    .S(_07419_),
    .Z(net248));
 MUX2_X1 _24778_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .B(net248),
    .S(_07420_),
    .Z(_01526_));
 MUX2_X1 _24779_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .B(_06818_),
    .S(_07419_),
    .Z(net249));
 MUX2_X1 _24780_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .B(net249),
    .S(_07420_),
    .Z(_01527_));
 MUX2_X1 _24781_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .B(_07124_),
    .S(_07419_),
    .Z(net250));
 MUX2_X1 _24782_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .B(net250),
    .S(_07420_),
    .Z(_01528_));
 MUX2_X1 _24783_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .B(_07126_),
    .S(_07419_),
    .Z(net251));
 MUX2_X1 _24784_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .B(net251),
    .S(_07420_),
    .Z(_01529_));
 MUX2_X1 _24785_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .B(_06828_),
    .S(_07419_),
    .Z(net252));
 MUX2_X1 _24786_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .B(net252),
    .S(_07420_),
    .Z(_01530_));
 MUX2_X1 _24787_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .B(_06839_),
    .S(_07419_),
    .Z(net253));
 MUX2_X1 _24788_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .B(net253),
    .S(_07420_),
    .Z(_01531_));
 NAND2_X1 _24789_ (.A1(_10319_),
    .A2(\load_store_unit_i.lsu_err_q ),
    .ZN(_07422_));
 NAND3_X1 _24790_ (.A1(_10324_),
    .A2(_10320_),
    .A3(_07422_),
    .ZN(_07423_));
 NAND3_X4 _24791_ (.A1(_10350_),
    .A2(_11427_),
    .A3(_06256_),
    .ZN(_07424_));
 NAND2_X1 _24792_ (.A1(_10320_),
    .A2(_03454_),
    .ZN(_07425_));
 NAND2_X1 _24793_ (.A1(_03453_),
    .A2(_10356_),
    .ZN(_07426_));
 OAI221_X1 _24794_ (.A(_07423_),
    .B1(_07424_),
    .B2(_07425_),
    .C1(net36),
    .C2(_07426_),
    .ZN(_07427_));
 INV_X1 _24795_ (.A(net37),
    .ZN(_07428_));
 NAND3_X1 _24796_ (.A1(_10322_),
    .A2(_03453_),
    .A3(_03454_),
    .ZN(_07429_));
 OAI21_X1 _24797_ (.A(_07428_),
    .B1(net36),
    .B2(_07429_),
    .ZN(_07430_));
 AND2_X1 _24798_ (.A1(_07427_),
    .A2(_07430_),
    .ZN(_07431_));
 CLKBUF_X2 _24799_ (.A(_07431_),
    .Z(_07432_));
 BUF_X4 _24800_ (.A(_07432_),
    .Z(_07433_));
 MUX2_X1 _24801_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .B(\alu_adder_result_ex[0] ),
    .S(_07433_),
    .Z(_01615_));
 MUX2_X1 _24802_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .B(net386),
    .S(_07433_),
    .Z(_01616_));
 MUX2_X1 _24803_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .B(\alu_adder_result_ex[11] ),
    .S(_07433_),
    .Z(_01617_));
 MUX2_X1 _24804_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .B(\alu_adder_result_ex[12] ),
    .S(_07433_),
    .Z(_01618_));
 MUX2_X1 _24805_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .B(\alu_adder_result_ex[13] ),
    .S(_07433_),
    .Z(_01619_));
 MUX2_X1 _24806_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .B(net380),
    .S(_07433_),
    .Z(_01620_));
 MUX2_X1 _24807_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .B(\alu_adder_result_ex[15] ),
    .S(_07433_),
    .Z(_01621_));
 MUX2_X1 _24808_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .B(\alu_adder_result_ex[16] ),
    .S(_07433_),
    .Z(_01622_));
 MUX2_X1 _24809_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .B(\alu_adder_result_ex[17] ),
    .S(_07433_),
    .Z(_01623_));
 MUX2_X1 _24810_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .B(net450),
    .S(_07433_),
    .Z(_01624_));
 CLKBUF_X3 _24811_ (.A(_07432_),
    .Z(_07434_));
 MUX2_X1 _24812_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .B(net381),
    .S(_07434_),
    .Z(_01625_));
 MUX2_X1 _24813_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .B(net15),
    .S(_07434_),
    .Z(_01626_));
 MUX2_X1 _24814_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .B(\alu_adder_result_ex[20] ),
    .S(_07434_),
    .Z(_01627_));
 MUX2_X1 _24815_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .B(net366),
    .S(_07434_),
    .Z(_01628_));
 MUX2_X1 _24816_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .B(\alu_adder_result_ex[22] ),
    .S(_07434_),
    .Z(_01629_));
 MUX2_X1 _24817_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .B(net372),
    .S(_07434_),
    .Z(_01630_));
 MUX2_X1 _24818_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .B(\alu_adder_result_ex[24] ),
    .S(_07434_),
    .Z(_01631_));
 MUX2_X1 _24819_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .B(net373),
    .S(_07434_),
    .Z(_01632_));
 MUX2_X1 _24820_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .B(net385),
    .S(_07434_),
    .Z(_01633_));
 MUX2_X1 _24821_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .B(\alu_adder_result_ex[27] ),
    .S(_07434_),
    .Z(_01634_));
 CLKBUF_X3 _24822_ (.A(_07432_),
    .Z(_07435_));
 MUX2_X1 _24823_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .B(\alu_adder_result_ex[28] ),
    .S(_07435_),
    .Z(_01635_));
 MUX2_X1 _24824_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .B(net14),
    .S(_07435_),
    .Z(_01636_));
 MUX2_X1 _24825_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .B(\alu_adder_result_ex[2] ),
    .S(_07435_),
    .Z(_01637_));
 MUX2_X1 _24826_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .B(\alu_adder_result_ex[30] ),
    .S(_07435_),
    .Z(_01638_));
 MUX2_X1 _24827_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .B(net279),
    .S(_07435_),
    .Z(_01639_));
 MUX2_X1 _24828_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .B(\alu_adder_result_ex[3] ),
    .S(_07435_),
    .Z(_01640_));
 MUX2_X1 _24829_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .B(\alu_adder_result_ex[4] ),
    .S(_07435_),
    .Z(_01641_));
 MUX2_X1 _24830_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .B(\alu_adder_result_ex[5] ),
    .S(_07435_),
    .Z(_01642_));
 MUX2_X1 _24831_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .B(\alu_adder_result_ex[6] ),
    .S(_07435_),
    .Z(_01643_));
 MUX2_X1 _24832_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .B(\alu_adder_result_ex[7] ),
    .S(_07435_),
    .Z(_01644_));
 MUX2_X1 _24833_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .B(\alu_adder_result_ex[8] ),
    .S(_07432_),
    .Z(_01645_));
 MUX2_X1 _24834_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .B(\alu_adder_result_ex[9] ),
    .S(_07432_),
    .Z(_01646_));
 NOR3_X1 _24835_ (.A1(_10287_),
    .A2(_10495_),
    .A3(_10909_),
    .ZN(_07436_));
 INV_X1 _24836_ (.A(_10320_),
    .ZN(_07437_));
 NOR2_X1 _24837_ (.A1(_07437_),
    .A2(_07428_),
    .ZN(_07438_));
 OAI21_X1 _24838_ (.A(_10325_),
    .B1(_10319_),
    .B2(_07424_),
    .ZN(_07439_));
 NAND2_X2 _24839_ (.A1(_07438_),
    .A2(_07439_),
    .ZN(_07440_));
 MUX2_X1 _24840_ (.A(_07436_),
    .B(\load_store_unit_i.data_sign_ext_q ),
    .S(_07440_),
    .Z(_01647_));
 NOR3_X4 _24841_ (.A1(_10289_),
    .A2(_10909_),
    .A3(_03434_),
    .ZN(net223));
 MUX2_X1 _24842_ (.A(net223),
    .B(\load_store_unit_i.data_we_q ),
    .S(_07440_),
    .Z(_01648_));
 AOI21_X4 _24843_ (.A(_07437_),
    .B1(_03454_),
    .B2(_07424_),
    .ZN(net190));
 INV_X1 _24844_ (.A(_10319_),
    .ZN(_07441_));
 NOR2_X1 _24845_ (.A1(_10324_),
    .A2(_07441_),
    .ZN(_07442_));
 AOI21_X1 _24846_ (.A(net37),
    .B1(_03453_),
    .B2(_07442_),
    .ZN(_07443_));
 INV_X1 _24847_ (.A(_07443_),
    .ZN(_07444_));
 AOI21_X1 _24848_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B1(net190),
    .B2(_07444_),
    .ZN(_07445_));
 CLKBUF_X2 _24849_ (.A(_16095_),
    .Z(_07446_));
 NOR2_X4 _24850_ (.A1(_10488_),
    .A2(_10909_),
    .ZN(_07447_));
 NAND3_X1 _24851_ (.A1(_10477_),
    .A2(_07446_),
    .A3(_07447_),
    .ZN(_07448_));
 OAI21_X2 _24852_ (.A(_07448_),
    .B1(_07447_),
    .B2(_03619_),
    .ZN(_07449_));
 OR2_X1 _24853_ (.A1(_10324_),
    .A2(_07449_),
    .ZN(_07450_));
 OAI21_X1 _24854_ (.A(_07441_),
    .B1(_07424_),
    .B2(_07450_),
    .ZN(_07451_));
 AOI21_X1 _24855_ (.A(_07445_),
    .B1(_07451_),
    .B2(_07438_),
    .ZN(_01649_));
 NAND2_X1 _24856_ (.A1(_10320_),
    .A2(_07428_),
    .ZN(_07452_));
 INV_X1 _24857_ (.A(_03453_),
    .ZN(_07453_));
 NAND3_X1 _24858_ (.A1(_10322_),
    .A2(_07453_),
    .A3(_03454_),
    .ZN(_07454_));
 AOI21_X1 _24859_ (.A(_10324_),
    .B1(_10319_),
    .B2(_07453_),
    .ZN(_07455_));
 OAI21_X1 _24860_ (.A(_07454_),
    .B1(_07455_),
    .B2(_07452_),
    .ZN(_07456_));
 AOI21_X2 _24861_ (.A(_07456_),
    .B1(_07424_),
    .B2(_03455_),
    .ZN(_07457_));
 OAI21_X1 _24862_ (.A(_07457_),
    .B1(_03453_),
    .B2(_07441_),
    .ZN(_07458_));
 AOI21_X1 _24863_ (.A(_07452_),
    .B1(_07458_),
    .B2(_10325_),
    .ZN(_01650_));
 AOI21_X1 _24864_ (.A(_10324_),
    .B1(net37),
    .B2(_07449_),
    .ZN(_07459_));
 NOR2_X1 _24865_ (.A1(_10319_),
    .A2(_07449_),
    .ZN(_07460_));
 AOI21_X1 _24866_ (.A(_07460_),
    .B1(_07442_),
    .B2(_03453_),
    .ZN(_07461_));
 OAI22_X1 _24867_ (.A1(_10319_),
    .A2(_07459_),
    .B1(_07461_),
    .B2(net37),
    .ZN(_07462_));
 NAND3_X1 _24868_ (.A1(_10320_),
    .A2(_07457_),
    .A3(_07462_),
    .ZN(_07463_));
 OAI21_X1 _24869_ (.A(_07463_),
    .B1(_07457_),
    .B2(_07441_),
    .ZN(_01651_));
 NOR3_X1 _24870_ (.A1(_10324_),
    .A2(_03453_),
    .A3(_10357_),
    .ZN(_07464_));
 MUX2_X1 _24871_ (.A(_10322_),
    .B(_07464_),
    .S(_07457_),
    .Z(_01652_));
 AOI21_X1 _24872_ (.A(_07426_),
    .B1(_07424_),
    .B2(_03455_),
    .ZN(_07465_));
 NAND2_X1 _24873_ (.A1(_03455_),
    .A2(_07424_),
    .ZN(_07466_));
 OAI21_X1 _24874_ (.A(_07426_),
    .B1(_07425_),
    .B2(_10322_),
    .ZN(_07467_));
 NAND2_X1 _24875_ (.A1(_07466_),
    .A2(_07467_),
    .ZN(_07468_));
 AOI22_X1 _24876_ (.A1(net36),
    .A2(_07465_),
    .B1(_07468_),
    .B2(\load_store_unit_i.lsu_err_q ),
    .ZN(_07469_));
 INV_X1 _24877_ (.A(_07469_),
    .ZN(_01653_));
 MUX2_X1 _24878_ (.A(\alu_adder_result_ex[0] ),
    .B(_04594_),
    .S(_07440_),
    .Z(_01654_));
 MUX2_X1 _24879_ (.A(net15),
    .B(_04597_),
    .S(_07440_),
    .Z(_01655_));
 OR2_X1 _24880_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_07426_),
    .ZN(_07470_));
 CLKBUF_X3 _24881_ (.A(_07470_),
    .Z(_07471_));
 BUF_X4 _24882_ (.A(_07471_),
    .Z(_07472_));
 MUX2_X1 _24883_ (.A(net67),
    .B(\load_store_unit_i.rdata_q[8] ),
    .S(_07472_),
    .Z(_01656_));
 MUX2_X1 _24884_ (.A(net47),
    .B(\load_store_unit_i.rdata_q[18] ),
    .S(_07472_),
    .Z(_01657_));
 MUX2_X1 _24885_ (.A(net48),
    .B(\load_store_unit_i.rdata_q[19] ),
    .S(_07472_),
    .Z(_01658_));
 MUX2_X1 _24886_ (.A(net50),
    .B(\load_store_unit_i.rdata_q[20] ),
    .S(_07472_),
    .Z(_01659_));
 MUX2_X1 _24887_ (.A(net51),
    .B(\load_store_unit_i.rdata_q[21] ),
    .S(_07472_),
    .Z(_01660_));
 MUX2_X1 _24888_ (.A(net52),
    .B(\load_store_unit_i.rdata_q[22] ),
    .S(_07472_),
    .Z(_01661_));
 MUX2_X1 _24889_ (.A(_04568_),
    .B(\load_store_unit_i.rdata_q[23] ),
    .S(_07472_),
    .Z(_01662_));
 MUX2_X1 _24890_ (.A(net53),
    .B(\load_store_unit_i.rdata_q[24] ),
    .S(_07472_),
    .Z(_01663_));
 MUX2_X1 _24891_ (.A(net54),
    .B(\load_store_unit_i.rdata_q[25] ),
    .S(_07472_),
    .Z(_01664_));
 MUX2_X1 _24892_ (.A(net55),
    .B(\load_store_unit_i.rdata_q[26] ),
    .S(_07472_),
    .Z(_01665_));
 BUF_X4 _24893_ (.A(_07471_),
    .Z(_07473_));
 MUX2_X1 _24894_ (.A(net56),
    .B(\load_store_unit_i.rdata_q[27] ),
    .S(_07473_),
    .Z(_01666_));
 MUX2_X1 _24895_ (.A(net68),
    .B(\load_store_unit_i.rdata_q[9] ),
    .S(_07473_),
    .Z(_01667_));
 MUX2_X1 _24896_ (.A(net57),
    .B(\load_store_unit_i.rdata_q[28] ),
    .S(_07473_),
    .Z(_01668_));
 MUX2_X1 _24897_ (.A(net58),
    .B(\load_store_unit_i.rdata_q[29] ),
    .S(_07473_),
    .Z(_01669_));
 MUX2_X1 _24898_ (.A(net60),
    .B(\load_store_unit_i.rdata_q[30] ),
    .S(_07473_),
    .Z(_01670_));
 MUX2_X1 _24899_ (.A(net61),
    .B(\load_store_unit_i.rdata_q[31] ),
    .S(_07473_),
    .Z(_01671_));
 MUX2_X1 _24900_ (.A(net39),
    .B(\load_store_unit_i.rdata_q[10] ),
    .S(_07473_),
    .Z(_01672_));
 MUX2_X1 _24901_ (.A(net40),
    .B(\load_store_unit_i.rdata_q[11] ),
    .S(_07473_),
    .Z(_01673_));
 MUX2_X1 _24902_ (.A(net41),
    .B(\load_store_unit_i.rdata_q[12] ),
    .S(_07473_),
    .Z(_01674_));
 MUX2_X1 _24903_ (.A(net42),
    .B(\load_store_unit_i.rdata_q[13] ),
    .S(_07473_),
    .Z(_01675_));
 MUX2_X1 _24904_ (.A(net43),
    .B(\load_store_unit_i.rdata_q[14] ),
    .S(_07471_),
    .Z(_01676_));
 MUX2_X1 _24905_ (.A(net44),
    .B(\load_store_unit_i.rdata_q[15] ),
    .S(_07471_),
    .Z(_01677_));
 MUX2_X1 _24906_ (.A(net45),
    .B(\load_store_unit_i.rdata_q[16] ),
    .S(_07471_),
    .Z(_01678_));
 MUX2_X1 _24907_ (.A(net46),
    .B(\load_store_unit_i.rdata_q[17] ),
    .S(_07471_),
    .Z(_01679_));
 NOR2_X1 _24908_ (.A1(_10909_),
    .A2(_10549_),
    .ZN(_07474_));
 MUX2_X1 _24909_ (.A(_07474_),
    .B(_04574_),
    .S(_07440_),
    .Z(_01680_));
 NOR2_X2 _24910_ (.A1(_10909_),
    .A2(_10677_),
    .ZN(_07475_));
 MUX2_X1 _24911_ (.A(_07475_),
    .B(_05270_),
    .S(_07440_),
    .Z(_01681_));
 MUX2_X1 _24912_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .S(_11429_),
    .Z(_01682_));
 MUX2_X1 _24913_ (.A(_11431_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_11429_),
    .Z(_01683_));
 MUX2_X1 _24914_ (.A(_06386_),
    .B(_03652_),
    .S(_03441_),
    .Z(_01684_));
 MUX2_X1 _24915_ (.A(_03617_),
    .B(_03611_),
    .S(_03441_),
    .Z(_01685_));
 MUX2_X1 _24916_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(_03647_),
    .S(_03441_),
    .Z(_01686_));
 BUF_X2 _24917_ (.A(_15530_),
    .Z(_07476_));
 CLKBUF_X2 _24918_ (.A(_07476_),
    .Z(_07477_));
 MUX2_X1 _24919_ (.A(_07477_),
    .B(_15526_),
    .S(_15842_),
    .Z(_07478_));
 BUF_X4 _24920_ (.A(_15524_),
    .Z(_07479_));
 BUF_X4 _24921_ (.A(_07479_),
    .Z(_07480_));
 BUF_X8 _24922_ (.A(_07480_),
    .Z(_07481_));
 OAI22_X4 _24923_ (.A1(_15842_),
    .A2(_05369_),
    .B1(_07478_),
    .B2(_07481_),
    .ZN(_07482_));
 INV_X1 _24924_ (.A(_07482_),
    .ZN(_07483_));
 OAI21_X2 _24925_ (.A(_03484_),
    .B1(_03507_),
    .B2(_04509_),
    .ZN(_07484_));
 OR2_X1 _24926_ (.A1(_15527_),
    .A2(_03486_),
    .ZN(_07485_));
 OR3_X1 _24927_ (.A1(_07484_),
    .A2(_03485_),
    .A3(_07485_),
    .ZN(_07486_));
 BUF_X4 _24928_ (.A(_07486_),
    .Z(_07487_));
 NOR2_X4 _24929_ (.A1(_04260_),
    .A2(_07487_),
    .ZN(_07488_));
 BUF_X8 _24930_ (.A(_07488_),
    .Z(_07489_));
 NAND2_X1 _24931_ (.A1(_05231_),
    .A2(_07489_),
    .ZN(_07490_));
 MUX2_X1 _24932_ (.A(_07483_),
    .B(\cs_registers_i.mcountinhibit[0] ),
    .S(_07490_),
    .Z(_01687_));
 MUX2_X1 _24933_ (.A(_15530_),
    .B(_11355_),
    .S(_15852_),
    .Z(_07491_));
 OAI22_X4 _24934_ (.A1(_15852_),
    .A2(_05461_),
    .B1(_07491_),
    .B2(_07479_),
    .ZN(_07492_));
 INV_X2 _24935_ (.A(_07492_),
    .ZN(_07493_));
 MUX2_X1 _24936_ (.A(_07493_),
    .B(\cs_registers_i.mcountinhibit[2] ),
    .S(_07490_),
    .Z(_01688_));
 NOR3_X2 _24937_ (.A1(_07484_),
    .A2(_03485_),
    .A3(_07485_),
    .ZN(_07494_));
 NAND4_X1 _24938_ (.A1(_03500_),
    .A2(_10922_),
    .A3(_11070_),
    .A4(_15873_),
    .ZN(_07495_));
 AOI21_X1 _24939_ (.A(_03499_),
    .B1(_15873_),
    .B2(_15857_),
    .ZN(_07496_));
 OAI21_X1 _24940_ (.A(_07495_),
    .B1(_07496_),
    .B2(_03500_),
    .ZN(_07497_));
 OAI21_X1 _24941_ (.A(_10922_),
    .B1(_03540_),
    .B2(_04289_),
    .ZN(_07498_));
 AND4_X1 _24942_ (.A1(_15509_),
    .A2(_15513_),
    .A3(_07497_),
    .A4(_07498_),
    .ZN(_07499_));
 NAND3_X1 _24943_ (.A1(_04237_),
    .A2(_07494_),
    .A3(_07499_),
    .ZN(_07500_));
 CLKBUF_X3 _24944_ (.A(_07500_),
    .Z(_07501_));
 CLKBUF_X3 _24945_ (.A(_07501_),
    .Z(_07502_));
 NAND2_X1 _24946_ (.A1(_00551_),
    .A2(_07502_),
    .ZN(_07503_));
 CLKBUF_X3 _24947_ (.A(_07501_),
    .Z(_07504_));
 OAI21_X1 _24948_ (.A(_07503_),
    .B1(_07504_),
    .B2(_07482_),
    .ZN(_07505_));
 MUX2_X1 _24949_ (.A(_04558_),
    .B(_00553_),
    .S(_07501_),
    .Z(_07506_));
 CLKBUF_X3 _24950_ (.A(_07506_),
    .Z(_07507_));
 MUX2_X1 _24951_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(_07505_),
    .S(_07507_),
    .Z(_01689_));
 MUX2_X2 _24952_ (.A(_05745_),
    .B(_05362_),
    .S(_07501_),
    .Z(_07508_));
 CLKBUF_X3 _24953_ (.A(_07508_),
    .Z(_07509_));
 INV_X1 _24954_ (.A(_05749_),
    .ZN(_07510_));
 NOR2_X4 _24955_ (.A1(_05748_),
    .A2(_05745_),
    .ZN(_07511_));
 NAND2_X2 _24956_ (.A1(_07494_),
    .A2(_07499_),
    .ZN(_07512_));
 NOR2_X2 _24957_ (.A1(_07511_),
    .A2(_07512_),
    .ZN(_07513_));
 CLKBUF_X2 _24958_ (.A(_15534_),
    .Z(_07514_));
 AND3_X1 _24959_ (.A1(_05459_),
    .A2(_05494_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .ZN(_07515_));
 NAND3_X2 _24960_ (.A1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .A2(_07514_),
    .A3(_07515_),
    .ZN(_07516_));
 INV_X1 _24961_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .ZN(_07517_));
 NAND3_X1 _24962_ (.A1(_05606_),
    .A2(_05628_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .ZN(_07518_));
 OR2_X1 _24963_ (.A1(_07517_),
    .A2(_07518_),
    .ZN(_07519_));
 OR2_X2 _24964_ (.A1(_07516_),
    .A2(_07519_),
    .ZN(_07520_));
 NOR3_X1 _24965_ (.A1(_07510_),
    .A2(_07513_),
    .A3(_07520_),
    .ZN(_07521_));
 NAND2_X1 _24966_ (.A1(_15921_),
    .A2(_05753_),
    .ZN(_07522_));
 MUX2_X1 _24967_ (.A(_15526_),
    .B(_07477_),
    .S(_15921_),
    .Z(_07523_));
 OAI21_X4 _24968_ (.A(_07522_),
    .B1(_07523_),
    .B2(_07481_),
    .ZN(_07524_));
 BUF_X4 _24969_ (.A(_07524_),
    .Z(_07525_));
 CLKBUF_X3 _24970_ (.A(_07513_),
    .Z(_07526_));
 AOI21_X1 _24971_ (.A(_07521_),
    .B1(_07525_),
    .B2(_07526_),
    .ZN(_07527_));
 CLKBUF_X3 _24972_ (.A(_07501_),
    .Z(_07528_));
 AOI21_X1 _24973_ (.A(_07508_),
    .B1(_07520_),
    .B2(_07528_),
    .ZN(_07529_));
 OAI22_X1 _24974_ (.A1(_07509_),
    .A2(_07527_),
    .B1(_07529_),
    .B2(_05749_),
    .ZN(_07530_));
 INV_X1 _24975_ (.A(_07530_),
    .ZN(_01690_));
 CLKBUF_X3 _24976_ (.A(_07513_),
    .Z(_07531_));
 CLKBUF_X2 _24977_ (.A(_11355_),
    .Z(_07532_));
 MUX2_X1 _24978_ (.A(_07532_),
    .B(_07476_),
    .S(_15928_),
    .Z(_07533_));
 BUF_X8 _24979_ (.A(_07479_),
    .Z(_07534_));
 OAI22_X4 _24980_ (.A1(_15924_),
    .A2(_05792_),
    .B1(_07533_),
    .B2(_07534_),
    .ZN(_07535_));
 NAND2_X1 _24981_ (.A1(_07531_),
    .A2(_07535_),
    .ZN(_07536_));
 CLKBUF_X3 _24982_ (.A(_07513_),
    .Z(_07537_));
 INV_X1 _24983_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .ZN(_07538_));
 NAND4_X2 _24984_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_05459_),
    .A3(_05494_),
    .A4(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .ZN(_07539_));
 NOR2_X1 _24985_ (.A1(_07538_),
    .A2(_07539_),
    .ZN(_07540_));
 NAND2_X2 _24986_ (.A1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .A2(_07540_),
    .ZN(_07541_));
 OR2_X2 _24987_ (.A1(_07519_),
    .A2(_07541_),
    .ZN(_07542_));
 NAND2_X1 _24988_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_05749_),
    .ZN(_07543_));
 OR3_X1 _24989_ (.A1(_07537_),
    .A2(_07542_),
    .A3(_07543_),
    .ZN(_07544_));
 AOI21_X1 _24990_ (.A(_07509_),
    .B1(_07536_),
    .B2(_07544_),
    .ZN(_07545_));
 CLKBUF_X3 _24991_ (.A(_07507_),
    .Z(_07546_));
 OAI21_X1 _24992_ (.A(_07504_),
    .B1(_07542_),
    .B2(_07510_),
    .ZN(_07547_));
 AOI21_X1 _24993_ (.A(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .B1(_07546_),
    .B2(_07547_),
    .ZN(_07548_));
 NOR2_X1 _24994_ (.A1(_07545_),
    .A2(_07548_),
    .ZN(_01691_));
 CLKBUF_X3 _24995_ (.A(_07506_),
    .Z(_07549_));
 CLKBUF_X3 _24996_ (.A(_07501_),
    .Z(_07550_));
 OAI21_X1 _24997_ (.A(_07550_),
    .B1(_07520_),
    .B2(_07543_),
    .ZN(_07551_));
 AOI21_X1 _24998_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B1(_07549_),
    .B2(_07551_),
    .ZN(_07552_));
 MUX2_X1 _24999_ (.A(_07532_),
    .B(_07476_),
    .S(_15936_),
    .Z(_07553_));
 OAI22_X4 _25000_ (.A1(_15932_),
    .A2(_05846_),
    .B1(_07553_),
    .B2(_07534_),
    .ZN(_07554_));
 NAND2_X1 _25001_ (.A1(_07526_),
    .A2(_07554_),
    .ZN(_07555_));
 NAND3_X2 _25002_ (.A1(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A3(_05749_),
    .ZN(_07556_));
 OR2_X1 _25003_ (.A1(_07537_),
    .A2(_07520_),
    .ZN(_07557_));
 OAI21_X1 _25004_ (.A(_07555_),
    .B1(_07556_),
    .B2(_07557_),
    .ZN(_07558_));
 CLKBUF_X3 _25005_ (.A(_07507_),
    .Z(_07559_));
 AOI21_X1 _25006_ (.A(_07552_),
    .B1(_07558_),
    .B2(_07559_),
    .ZN(_01692_));
 CLKBUF_X3 _25007_ (.A(_07507_),
    .Z(_07560_));
 OAI21_X1 _25008_ (.A(_07528_),
    .B1(_07542_),
    .B2(_07556_),
    .ZN(_07561_));
 AOI21_X1 _25009_ (.A(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .B1(_07560_),
    .B2(_07561_),
    .ZN(_07562_));
 CLKBUF_X3 _25010_ (.A(_07501_),
    .Z(_07563_));
 CLKBUF_X2 _25011_ (.A(_15530_),
    .Z(_07564_));
 MUX2_X1 _25012_ (.A(_11356_),
    .B(_07564_),
    .S(_15944_),
    .Z(_07565_));
 NOR2_X1 _25013_ (.A1(_07480_),
    .A2(_07565_),
    .ZN(_07566_));
 NOR3_X2 _25014_ (.A1(_05877_),
    .A2(_05880_),
    .A3(_05886_),
    .ZN(_07567_));
 AOI21_X2 _25015_ (.A(_07566_),
    .B1(_07567_),
    .B2(_15944_),
    .ZN(_07568_));
 BUF_X4 _25016_ (.A(_07568_),
    .Z(_07569_));
 OR2_X1 _25017_ (.A1(_07563_),
    .A2(_07569_),
    .ZN(_07570_));
 INV_X1 _25018_ (.A(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .ZN(_07571_));
 OR4_X1 _25019_ (.A1(_07571_),
    .A2(_07513_),
    .A3(_07542_),
    .A4(_07556_),
    .ZN(_07572_));
 AOI21_X1 _25020_ (.A(_07509_),
    .B1(_07570_),
    .B2(_07572_),
    .ZN(_07573_));
 NOR2_X1 _25021_ (.A1(_07562_),
    .A2(_07573_),
    .ZN(_01693_));
 NAND4_X2 _25022_ (.A1(_15509_),
    .A2(_15513_),
    .A3(_07497_),
    .A4(_07498_),
    .ZN(_07574_));
 OAI33_X1 _25023_ (.A1(_07511_),
    .A2(_07487_),
    .A3(_07574_),
    .B1(_07520_),
    .B2(_07556_),
    .B3(_07571_),
    .ZN(_07575_));
 AOI21_X1 _25024_ (.A(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .B1(_07549_),
    .B2(_07575_),
    .ZN(_07576_));
 MUX2_X1 _25025_ (.A(_11356_),
    .B(_07476_),
    .S(_15952_),
    .Z(_07577_));
 NOR2_X1 _25026_ (.A1(_07534_),
    .A2(_07577_),
    .ZN(_07578_));
 AOI21_X4 _25027_ (.A(_07578_),
    .B1(_05924_),
    .B2(_15952_),
    .ZN(_07579_));
 OR2_X1 _25028_ (.A1(_07563_),
    .A2(_07579_),
    .ZN(_07580_));
 NOR2_X1 _25029_ (.A1(_07571_),
    .A2(_07556_),
    .ZN(_07581_));
 NAND2_X1 _25030_ (.A1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .A2(_07581_),
    .ZN(_07582_));
 OAI21_X1 _25031_ (.A(_07580_),
    .B1(_07582_),
    .B2(_07557_),
    .ZN(_07583_));
 AOI21_X1 _25032_ (.A(_07576_),
    .B1(_07583_),
    .B2(_07559_),
    .ZN(_01694_));
 MUX2_X1 _25033_ (.A(_11356_),
    .B(_07564_),
    .S(_15957_),
    .Z(_07584_));
 OAI22_X4 _25034_ (.A1(_15961_),
    .A2(_05970_),
    .B1(_07584_),
    .B2(_07480_),
    .ZN(_07585_));
 NAND2_X1 _25035_ (.A1(_07537_),
    .A2(_07585_),
    .ZN(_07586_));
 NOR2_X1 _25036_ (.A1(_07542_),
    .A2(_07582_),
    .ZN(_07587_));
 NAND3_X1 _25037_ (.A1(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .A2(_07550_),
    .A3(_07587_),
    .ZN(_07588_));
 AOI21_X1 _25038_ (.A(_07509_),
    .B1(_07586_),
    .B2(_07588_),
    .ZN(_07589_));
 CLKBUF_X3 _25039_ (.A(_07537_),
    .Z(_07590_));
 OAI21_X1 _25040_ (.A(_07546_),
    .B1(_07587_),
    .B2(_07590_),
    .ZN(_07591_));
 INV_X1 _25041_ (.A(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .ZN(_07592_));
 AOI21_X1 _25042_ (.A(_07589_),
    .B1(_07591_),
    .B2(_07592_),
    .ZN(_01695_));
 INV_X1 _25043_ (.A(_06004_),
    .ZN(_07593_));
 NAND3_X2 _25044_ (.A1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .A3(_07581_),
    .ZN(_07594_));
 NOR2_X1 _25045_ (.A1(_07520_),
    .A2(_07594_),
    .ZN(_07595_));
 CLKBUF_X3 _25046_ (.A(_07537_),
    .Z(_07596_));
 OAI21_X1 _25047_ (.A(_07546_),
    .B1(_07595_),
    .B2(_07596_),
    .ZN(_07597_));
 MUX2_X1 _25048_ (.A(_11356_),
    .B(_07564_),
    .S(_15968_),
    .Z(_07598_));
 NOR2_X1 _25049_ (.A1(_07534_),
    .A2(_07598_),
    .ZN(_07599_));
 AOI21_X4 _25050_ (.A(_07599_),
    .B1(_06013_),
    .B2(_15968_),
    .ZN(_07600_));
 OR2_X1 _25051_ (.A1(_07563_),
    .A2(_07600_),
    .ZN(_07601_));
 NAND2_X1 _25052_ (.A1(_06004_),
    .A2(_07595_),
    .ZN(_07602_));
 OAI21_X1 _25053_ (.A(_07601_),
    .B1(_07602_),
    .B2(_07596_),
    .ZN(_07603_));
 AOI22_X1 _25054_ (.A1(_07593_),
    .A2(_07597_),
    .B1(_07603_),
    .B2(_07560_),
    .ZN(_01696_));
 MUX2_X1 _25055_ (.A(_07532_),
    .B(_07476_),
    .S(_15976_),
    .Z(_07604_));
 OAI22_X4 _25056_ (.A1(_15972_),
    .A2(_06054_),
    .B1(_07604_),
    .B2(_07534_),
    .ZN(_07605_));
 NAND2_X1 _25057_ (.A1(_07531_),
    .A2(_07605_),
    .ZN(_07606_));
 NOR3_X1 _25058_ (.A1(_07593_),
    .A2(_07542_),
    .A3(_07594_),
    .ZN(_07607_));
 NAND3_X1 _25059_ (.A1(_06037_),
    .A2(_07550_),
    .A3(_07607_),
    .ZN(_07608_));
 AOI21_X1 _25060_ (.A(_07508_),
    .B1(_07606_),
    .B2(_07608_),
    .ZN(_07609_));
 OAI21_X1 _25061_ (.A(_07546_),
    .B1(_07607_),
    .B2(_07590_),
    .ZN(_07610_));
 INV_X1 _25062_ (.A(_06037_),
    .ZN(_07611_));
 AOI21_X1 _25063_ (.A(_07609_),
    .B1(_07610_),
    .B2(_07611_),
    .ZN(_01697_));
 OAI21_X1 _25064_ (.A(_07550_),
    .B1(_07602_),
    .B2(_07611_),
    .ZN(_07612_));
 AOI21_X1 _25065_ (.A(_06094_),
    .B1(_07549_),
    .B2(_07612_),
    .ZN(_07613_));
 AND4_X1 _25066_ (.A1(_06004_),
    .A2(_06037_),
    .A3(_06094_),
    .A4(_07595_),
    .ZN(_07614_));
 MUX2_X1 _25067_ (.A(_11356_),
    .B(_07564_),
    .S(_15981_),
    .Z(_07615_));
 OAI22_X4 _25068_ (.A1(_15985_),
    .A2(_06097_),
    .B1(_07615_),
    .B2(_07479_),
    .ZN(_07616_));
 AND2_X1 _25069_ (.A1(_04756_),
    .A2(_03532_),
    .ZN(_07617_));
 NAND2_X1 _25070_ (.A1(_03518_),
    .A2(_11427_),
    .ZN(_07618_));
 OR4_X2 _25071_ (.A1(_15527_),
    .A2(_07484_),
    .A3(_03485_),
    .A4(_07618_),
    .ZN(_07619_));
 NOR3_X2 _25072_ (.A1(_07617_),
    .A2(_07619_),
    .A3(_07574_),
    .ZN(_07620_));
 MUX2_X1 _25073_ (.A(_07614_),
    .B(_07616_),
    .S(_07620_),
    .Z(_07621_));
 AOI21_X1 _25074_ (.A(_07613_),
    .B1(_07621_),
    .B2(_07559_),
    .ZN(_01698_));
 MUX2_X1 _25075_ (.A(_07532_),
    .B(_07477_),
    .S(_15992_),
    .Z(_07622_));
 OAI22_X4 _25076_ (.A1(_15988_),
    .A2(_06127_),
    .B1(_07622_),
    .B2(_07481_),
    .ZN(_07623_));
 BUF_X4 _25077_ (.A(_07623_),
    .Z(_07624_));
 NAND2_X1 _25078_ (.A1(_07531_),
    .A2(_07624_),
    .ZN(_07625_));
 NOR2_X1 _25079_ (.A1(_07542_),
    .A2(_07594_),
    .ZN(_07626_));
 AND4_X2 _25080_ (.A1(_06004_),
    .A2(_06037_),
    .A3(_06094_),
    .A4(_07626_),
    .ZN(_07627_));
 NAND2_X1 _25081_ (.A1(_07502_),
    .A2(_07627_),
    .ZN(_07628_));
 INV_X1 _25082_ (.A(_06123_),
    .ZN(_07629_));
 OAI21_X1 _25083_ (.A(_07625_),
    .B1(_07628_),
    .B2(_07629_),
    .ZN(_07630_));
 OAI21_X1 _25084_ (.A(_07507_),
    .B1(_07627_),
    .B2(_07596_),
    .ZN(_07631_));
 AOI22_X1 _25085_ (.A1(_07559_),
    .A2(_07630_),
    .B1(_07631_),
    .B2(_07629_),
    .ZN(_01699_));
 NAND2_X1 _25086_ (.A1(_15535_),
    .A2(_07563_),
    .ZN(_07632_));
 MUX2_X1 _25087_ (.A(_07477_),
    .B(_15526_),
    .S(_15845_),
    .Z(_07633_));
 OAI22_X2 _25088_ (.A1(_15845_),
    .A2(_05407_),
    .B1(_07633_),
    .B2(_07481_),
    .ZN(_07634_));
 BUF_X4 _25089_ (.A(_07634_),
    .Z(_07635_));
 CLKBUF_X3 _25090_ (.A(_07501_),
    .Z(_07636_));
 OAI21_X1 _25091_ (.A(_07632_),
    .B1(_07635_),
    .B2(_07636_),
    .ZN(_07637_));
 MUX2_X1 _25092_ (.A(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .B(_07637_),
    .S(_07507_),
    .Z(_01700_));
 MUX2_X1 _25093_ (.A(_07532_),
    .B(_07476_),
    .S(_15997_),
    .Z(_07638_));
 OAI22_X4 _25094_ (.A1(_16001_),
    .A2(_06170_),
    .B1(_07638_),
    .B2(_07534_),
    .ZN(_07639_));
 BUF_X4 _25095_ (.A(_07639_),
    .Z(_07640_));
 NAND2_X1 _25096_ (.A1(_07526_),
    .A2(_07640_),
    .ZN(_07641_));
 NAND4_X1 _25097_ (.A1(_06123_),
    .A2(_06168_),
    .A3(_07636_),
    .A4(_07614_),
    .ZN(_07642_));
 AOI21_X1 _25098_ (.A(_07509_),
    .B1(_07641_),
    .B2(_07642_),
    .ZN(_07643_));
 INV_X1 _25099_ (.A(_07614_),
    .ZN(_07644_));
 OAI21_X1 _25100_ (.A(_07504_),
    .B1(_07644_),
    .B2(_07629_),
    .ZN(_07645_));
 AOI21_X1 _25101_ (.A(_06168_),
    .B1(_07546_),
    .B2(_07645_),
    .ZN(_07646_));
 NOR2_X1 _25102_ (.A1(_07643_),
    .A2(_07646_),
    .ZN(_01701_));
 NAND3_X1 _25103_ (.A1(_06123_),
    .A2(_06168_),
    .A3(_07627_),
    .ZN(_07647_));
 NAND2_X1 _25104_ (.A1(_07504_),
    .A2(_07647_),
    .ZN(_07648_));
 AOI21_X1 _25105_ (.A(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .B1(_07549_),
    .B2(_07648_),
    .ZN(_07649_));
 MUX2_X1 _25106_ (.A(_11355_),
    .B(_07564_),
    .S(_16005_),
    .Z(_07650_));
 OAI22_X4 _25107_ (.A1(_16009_),
    .A2(_06197_),
    .B1(_07650_),
    .B2(_07479_),
    .ZN(_07651_));
 NAND2_X1 _25108_ (.A1(_07537_),
    .A2(_07651_),
    .ZN(_07652_));
 NAND3_X2 _25109_ (.A1(_06123_),
    .A2(_06168_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .ZN(_07653_));
 OAI21_X1 _25110_ (.A(_07652_),
    .B1(_07653_),
    .B2(_07628_),
    .ZN(_07654_));
 AOI21_X1 _25111_ (.A(_07649_),
    .B1(_07654_),
    .B2(_07559_),
    .ZN(_01702_));
 MUX2_X1 _25112_ (.A(_07476_),
    .B(_07532_),
    .S(_16017_),
    .Z(_07655_));
 OAI22_X4 _25113_ (.A1(_16017_),
    .A2(_04562_),
    .B1(_07655_),
    .B2(_07534_),
    .ZN(_07656_));
 BUF_X4 _25114_ (.A(_07656_),
    .Z(_07657_));
 NAND2_X1 _25115_ (.A1(_07537_),
    .A2(_07657_),
    .ZN(_07658_));
 INV_X1 _25116_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .ZN(_07659_));
 NOR2_X2 _25117_ (.A1(_07659_),
    .A2(_07653_),
    .ZN(_07660_));
 NAND3_X1 _25118_ (.A1(_07528_),
    .A2(_07614_),
    .A3(_07660_),
    .ZN(_07661_));
 AOI21_X1 _25119_ (.A(_07509_),
    .B1(_07658_),
    .B2(_07661_),
    .ZN(_07662_));
 OAI21_X1 _25120_ (.A(_07504_),
    .B1(_07644_),
    .B2(_07653_),
    .ZN(_07663_));
 AOI21_X1 _25121_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B1(_07546_),
    .B2(_07663_),
    .ZN(_07664_));
 NOR2_X1 _25122_ (.A1(_07662_),
    .A2(_07664_),
    .ZN(_01703_));
 NAND2_X1 _25123_ (.A1(_07627_),
    .A2(_07660_),
    .ZN(_07665_));
 NAND2_X1 _25124_ (.A1(_07504_),
    .A2(_07665_),
    .ZN(_07666_));
 AOI21_X1 _25125_ (.A(_04758_),
    .B1(_07549_),
    .B2(_07666_),
    .ZN(_07667_));
 MUX2_X1 _25126_ (.A(_07564_),
    .B(_11356_),
    .S(_16020_),
    .Z(_07668_));
 OAI22_X4 _25127_ (.A1(_16020_),
    .A2(_04762_),
    .B1(_07668_),
    .B2(_07480_),
    .ZN(_07669_));
 NAND2_X1 _25128_ (.A1(_07531_),
    .A2(_07669_),
    .ZN(_07670_));
 NAND2_X1 _25129_ (.A1(_04758_),
    .A2(_07660_),
    .ZN(_07671_));
 OAI21_X1 _25130_ (.A(_07670_),
    .B1(_07671_),
    .B2(_07628_),
    .ZN(_07672_));
 AOI21_X1 _25131_ (.A(_07667_),
    .B1(_07672_),
    .B2(_07559_),
    .ZN(_01704_));
 OAI21_X1 _25132_ (.A(_07550_),
    .B1(_07644_),
    .B2(_07671_),
    .ZN(_07673_));
 AOI21_X1 _25133_ (.A(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .B1(_07549_),
    .B2(_07673_),
    .ZN(_07674_));
 MUX2_X1 _25134_ (.A(_07564_),
    .B(_11356_),
    .S(_16033_),
    .Z(_07675_));
 OAI22_X4 _25135_ (.A1(_16033_),
    .A2(_04903_),
    .B1(_07675_),
    .B2(_07480_),
    .ZN(_07676_));
 NAND2_X1 _25136_ (.A1(_07531_),
    .A2(_07676_),
    .ZN(_07677_));
 NAND4_X1 _25137_ (.A1(_04758_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A3(_07614_),
    .A4(_07660_),
    .ZN(_07678_));
 OAI21_X1 _25138_ (.A(_07677_),
    .B1(_07678_),
    .B2(_07590_),
    .ZN(_07679_));
 AOI21_X1 _25139_ (.A(_07674_),
    .B1(_07679_),
    .B2(_07559_),
    .ZN(_01705_));
 CLKBUF_X3 _25140_ (.A(_07501_),
    .Z(_07680_));
 INV_X1 _25141_ (.A(_07627_),
    .ZN(_07681_));
 NAND3_X2 _25142_ (.A1(_04758_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A3(_07660_),
    .ZN(_07682_));
 OAI21_X1 _25143_ (.A(_07680_),
    .B1(_07681_),
    .B2(_07682_),
    .ZN(_07683_));
 AOI21_X1 _25144_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .B1(_07549_),
    .B2(_07683_),
    .ZN(_07684_));
 MUX2_X1 _25145_ (.A(_11355_),
    .B(_15530_),
    .S(_16040_),
    .Z(_07685_));
 NOR2_X1 _25146_ (.A1(_07480_),
    .A2(_07685_),
    .ZN(_07686_));
 NOR3_X4 _25147_ (.A1(_04962_),
    .A2(_04966_),
    .A3(_04974_),
    .ZN(_07687_));
 AOI21_X4 _25148_ (.A(_07686_),
    .B1(_07687_),
    .B2(_16040_),
    .ZN(_07688_));
 BUF_X4 _25149_ (.A(_07688_),
    .Z(_07689_));
 OR2_X1 _25150_ (.A1(_07563_),
    .A2(_07689_),
    .ZN(_07690_));
 NAND4_X2 _25151_ (.A1(_06004_),
    .A2(_06037_),
    .A3(_06094_),
    .A4(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .ZN(_07691_));
 OR4_X2 _25152_ (.A1(_07519_),
    .A2(_07594_),
    .A3(_07682_),
    .A4(_07691_),
    .ZN(_07692_));
 OR2_X2 _25153_ (.A1(_07541_),
    .A2(_07692_),
    .ZN(_07693_));
 OAI21_X1 _25154_ (.A(_07690_),
    .B1(_07693_),
    .B2(_07590_),
    .ZN(_07694_));
 AOI21_X1 _25155_ (.A(_07684_),
    .B1(_07694_),
    .B2(_07559_),
    .ZN(_01706_));
 MUX2_X1 _25156_ (.A(_15526_),
    .B(_07477_),
    .S(_16045_),
    .Z(_07695_));
 OAI22_X4 _25157_ (.A1(_16049_),
    .A2(_05034_),
    .B1(_07695_),
    .B2(_07481_),
    .ZN(_07696_));
 NAND2_X1 _25158_ (.A1(_07537_),
    .A2(_07696_),
    .ZN(_07697_));
 NOR2_X2 _25159_ (.A1(_07516_),
    .A2(_07692_),
    .ZN(_07698_));
 NAND3_X1 _25160_ (.A1(_05032_),
    .A2(_07550_),
    .A3(_07698_),
    .ZN(_07699_));
 AOI21_X1 _25161_ (.A(_07508_),
    .B1(_07697_),
    .B2(_07699_),
    .ZN(_07700_));
 OAI21_X1 _25162_ (.A(_07546_),
    .B1(_07698_),
    .B2(_07590_),
    .ZN(_07701_));
 INV_X1 _25163_ (.A(_05032_),
    .ZN(_07702_));
 AOI21_X1 _25164_ (.A(_07700_),
    .B1(_07701_),
    .B2(_07702_),
    .ZN(_01707_));
 OAI33_X1 _25165_ (.A1(_07617_),
    .A2(_07619_),
    .A3(_07574_),
    .B1(_07541_),
    .B2(_07692_),
    .B3(_07702_),
    .ZN(_07703_));
 AOI21_X1 _25166_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B1(_07549_),
    .B2(_07703_),
    .ZN(_07704_));
 NAND2_X2 _25167_ (.A1(_05032_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .ZN(_07705_));
 NOR2_X1 _25168_ (.A1(_07693_),
    .A2(_07705_),
    .ZN(_07706_));
 MUX2_X1 _25169_ (.A(_07532_),
    .B(_07476_),
    .S(_16056_),
    .Z(_07707_));
 OAI22_X4 _25170_ (.A1(_16052_),
    .A2(_04787_),
    .B1(_07707_),
    .B2(_07534_),
    .ZN(_07708_));
 BUF_X4 _25171_ (.A(_07708_),
    .Z(_07709_));
 MUX2_X1 _25172_ (.A(_07706_),
    .B(_07709_),
    .S(_07620_),
    .Z(_07710_));
 AOI21_X1 _25173_ (.A(_07704_),
    .B1(_07710_),
    .B2(_07560_),
    .ZN(_01708_));
 CLKBUF_X3 _25174_ (.A(_07563_),
    .Z(_07711_));
 NAND3_X2 _25175_ (.A1(_05032_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .A3(_07698_),
    .ZN(_07712_));
 NAND2_X1 _25176_ (.A1(_07711_),
    .A2(_07712_),
    .ZN(_07713_));
 AOI21_X1 _25177_ (.A(_05066_),
    .B1(_07560_),
    .B2(_07713_),
    .ZN(_07714_));
 MUX2_X1 _25178_ (.A(_15530_),
    .B(_11355_),
    .S(_16060_),
    .Z(_07715_));
 NOR2_X1 _25179_ (.A1(_07480_),
    .A2(_07715_),
    .ZN(_07716_));
 AOI21_X2 _25180_ (.A(_07716_),
    .B1(_05077_),
    .B2(_16064_),
    .ZN(_07717_));
 BUF_X4 _25181_ (.A(_07717_),
    .Z(_07718_));
 OR2_X1 _25182_ (.A1(_07563_),
    .A2(_07718_),
    .ZN(_07719_));
 INV_X1 _25183_ (.A(_07712_),
    .ZN(_07720_));
 NAND3_X1 _25184_ (.A1(_05066_),
    .A2(_07504_),
    .A3(_07720_),
    .ZN(_07721_));
 AOI21_X1 _25185_ (.A(_07509_),
    .B1(_07719_),
    .B2(_07721_),
    .ZN(_07722_));
 NOR2_X1 _25186_ (.A1(_07714_),
    .A2(_07722_),
    .ZN(_01709_));
 NAND2_X1 _25187_ (.A1(_05066_),
    .A2(_07706_),
    .ZN(_07723_));
 NAND2_X1 _25188_ (.A1(_07711_),
    .A2(_07723_),
    .ZN(_07724_));
 AOI21_X1 _25189_ (.A(_05142_),
    .B1(_07560_),
    .B2(_07724_),
    .ZN(_07725_));
 MUX2_X1 _25190_ (.A(_07477_),
    .B(_07532_),
    .S(_16068_),
    .Z(_07726_));
 OAI22_X4 _25191_ (.A1(_16068_),
    .A2(_05145_),
    .B1(_07726_),
    .B2(_07481_),
    .ZN(_07727_));
 BUF_X4 _25192_ (.A(_07727_),
    .Z(_07728_));
 NAND2_X1 _25193_ (.A1(_07526_),
    .A2(_07728_),
    .ZN(_07729_));
 NAND4_X1 _25194_ (.A1(_05066_),
    .A2(_05142_),
    .A3(_07550_),
    .A4(_07706_),
    .ZN(_07730_));
 AOI21_X1 _25195_ (.A(_07509_),
    .B1(_07729_),
    .B2(_07730_),
    .ZN(_07731_));
 NOR2_X1 _25196_ (.A1(_07725_),
    .A2(_07731_),
    .ZN(_01710_));
 NAND2_X1 _25197_ (.A1(_07492_),
    .A2(_07537_),
    .ZN(_07732_));
 NAND3_X1 _25198_ (.A1(_05459_),
    .A2(_07514_),
    .A3(_07502_),
    .ZN(_07733_));
 AOI21_X1 _25199_ (.A(_07508_),
    .B1(_07732_),
    .B2(_07733_),
    .ZN(_07734_));
 OAI21_X1 _25200_ (.A(_07546_),
    .B1(_07590_),
    .B2(_07514_),
    .ZN(_07735_));
 INV_X1 _25201_ (.A(_05459_),
    .ZN(_07736_));
 AOI21_X1 _25202_ (.A(_07734_),
    .B1(_07735_),
    .B2(_07736_),
    .ZN(_01711_));
 CLKBUF_X3 _25203_ (.A(_07501_),
    .Z(_07737_));
 NAND3_X1 _25204_ (.A1(_05066_),
    .A2(_05142_),
    .A3(_07720_),
    .ZN(_07738_));
 NAND2_X1 _25205_ (.A1(_07737_),
    .A2(_07738_),
    .ZN(_07739_));
 AOI21_X1 _25206_ (.A(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .B1(_07549_),
    .B2(_07739_),
    .ZN(_07740_));
 NAND3_X4 _25207_ (.A1(_05066_),
    .A2(_05142_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .ZN(_07741_));
 NOR2_X2 _25208_ (.A1(_07712_),
    .A2(_07741_),
    .ZN(_07742_));
 NAND2_X1 _25209_ (.A1(_16080_),
    .A2(_05203_),
    .ZN(_07743_));
 MUX2_X1 _25210_ (.A(_15526_),
    .B(_07477_),
    .S(_16080_),
    .Z(_07744_));
 OAI21_X4 _25211_ (.A(_07743_),
    .B1(_07744_),
    .B2(_07481_),
    .ZN(_07745_));
 MUX2_X1 _25212_ (.A(_07742_),
    .B(_07745_),
    .S(_07620_),
    .Z(_07746_));
 AOI21_X1 _25213_ (.A(_07740_),
    .B1(_07746_),
    .B2(_07560_),
    .ZN(_01712_));
 MUX2_X1 _25214_ (.A(_07476_),
    .B(_07532_),
    .S(_15496_),
    .Z(_07747_));
 OAI22_X4 _25215_ (.A1(_15496_),
    .A2(_05238_),
    .B1(_07747_),
    .B2(_07534_),
    .ZN(_07748_));
 NAND2_X1 _25216_ (.A1(_07531_),
    .A2(_07748_),
    .ZN(_07749_));
 NOR3_X4 _25217_ (.A1(_07693_),
    .A2(_07705_),
    .A3(_07741_),
    .ZN(_07750_));
 NAND3_X1 _25218_ (.A1(_05236_),
    .A2(_07550_),
    .A3(_07750_),
    .ZN(_07751_));
 AOI21_X1 _25219_ (.A(_07508_),
    .B1(_07749_),
    .B2(_07751_),
    .ZN(_07752_));
 OAI21_X1 _25220_ (.A(_07546_),
    .B1(_07750_),
    .B2(_07590_),
    .ZN(_07753_));
 INV_X1 _25221_ (.A(_05236_),
    .ZN(_07754_));
 AOI21_X1 _25222_ (.A(_07752_),
    .B1(_07753_),
    .B2(_07754_),
    .ZN(_01713_));
 OAI21_X1 _25223_ (.A(_00553_),
    .B1(_04560_),
    .B2(_07512_),
    .ZN(_07755_));
 OAI21_X2 _25224_ (.A(_07755_),
    .B1(_07512_),
    .B2(_04558_),
    .ZN(_07756_));
 BUF_X2 _25225_ (.A(_07756_),
    .Z(_07757_));
 CLKBUF_X3 _25226_ (.A(_07757_),
    .Z(_07758_));
 NAND2_X1 _25227_ (.A1(_05236_),
    .A2(_07742_),
    .ZN(_07759_));
 NAND2_X1 _25228_ (.A1(_07711_),
    .A2(_07759_),
    .ZN(_07760_));
 AOI21_X1 _25229_ (.A(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .B1(_07758_),
    .B2(_07760_),
    .ZN(_07761_));
 INV_X2 _25230_ (.A(_07756_),
    .ZN(_07762_));
 NAND2_X1 _25231_ (.A1(_07482_),
    .A2(_07526_),
    .ZN(_07763_));
 AND2_X2 _25232_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(_05236_),
    .ZN(_07764_));
 NAND3_X1 _25233_ (.A1(_07528_),
    .A2(_07742_),
    .A3(_07764_),
    .ZN(_07765_));
 AOI21_X1 _25234_ (.A(_07762_),
    .B1(_07763_),
    .B2(_07765_),
    .ZN(_07766_));
 NOR2_X1 _25235_ (.A1(_07761_),
    .A2(_07766_),
    .ZN(_01714_));
 CLKBUF_X3 _25236_ (.A(_07757_),
    .Z(_07767_));
 NAND2_X1 _25237_ (.A1(_07750_),
    .A2(_07764_),
    .ZN(_07768_));
 NAND2_X1 _25238_ (.A1(_07737_),
    .A2(_07768_),
    .ZN(_07769_));
 AOI21_X1 _25239_ (.A(_05404_),
    .B1(_07767_),
    .B2(_07769_),
    .ZN(_07770_));
 NAND2_X1 _25240_ (.A1(_07526_),
    .A2(_07635_),
    .ZN(_07771_));
 INV_X1 _25241_ (.A(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .ZN(_07772_));
 NOR3_X2 _25242_ (.A1(_07538_),
    .A2(_07772_),
    .A3(_07539_),
    .ZN(_07773_));
 NOR4_X2 _25243_ (.A1(_07519_),
    .A2(_07594_),
    .A3(_07682_),
    .A4(_07691_),
    .ZN(_07774_));
 NAND2_X1 _25244_ (.A1(_07773_),
    .A2(_07774_),
    .ZN(_07775_));
 NOR3_X2 _25245_ (.A1(_07775_),
    .A2(_07705_),
    .A3(_07741_),
    .ZN(_07776_));
 NAND3_X1 _25246_ (.A1(_05404_),
    .A2(_07776_),
    .A3(_07764_),
    .ZN(_07777_));
 OAI21_X1 _25247_ (.A(_07771_),
    .B1(_07777_),
    .B2(_07590_),
    .ZN(_07778_));
 CLKBUF_X3 _25248_ (.A(_07757_),
    .Z(_07779_));
 AOI21_X1 _25249_ (.A(_07770_),
    .B1(_07778_),
    .B2(_07779_),
    .ZN(_01715_));
 NAND3_X1 _25250_ (.A1(_05404_),
    .A2(_07742_),
    .A3(_07764_),
    .ZN(_07780_));
 NAND2_X1 _25251_ (.A1(_07711_),
    .A2(_07780_),
    .ZN(_07781_));
 AOI21_X1 _25252_ (.A(_05457_),
    .B1(_07758_),
    .B2(_07781_),
    .ZN(_07782_));
 INV_X1 _25253_ (.A(_05457_),
    .ZN(_07783_));
 NOR2_X2 _25254_ (.A1(_07783_),
    .A2(_07780_),
    .ZN(_07784_));
 NAND2_X1 _25255_ (.A1(_07528_),
    .A2(_07784_),
    .ZN(_07785_));
 AOI21_X1 _25256_ (.A(_07762_),
    .B1(_07785_),
    .B2(_07732_),
    .ZN(_07786_));
 NOR2_X1 _25257_ (.A1(_07782_),
    .A2(_07786_),
    .ZN(_01716_));
 NAND4_X2 _25258_ (.A1(_05404_),
    .A2(_05457_),
    .A3(_07750_),
    .A4(_07764_),
    .ZN(_07787_));
 NAND2_X1 _25259_ (.A1(_07737_),
    .A2(_07787_),
    .ZN(_07788_));
 AOI21_X1 _25260_ (.A(_05482_),
    .B1(_07767_),
    .B2(_07788_),
    .ZN(_07789_));
 MUX2_X1 _25261_ (.A(_07564_),
    .B(_11355_),
    .S(_15865_),
    .Z(_07790_));
 OAI22_X4 _25262_ (.A1(_15865_),
    .A2(_05497_),
    .B1(_07790_),
    .B2(_07480_),
    .ZN(_07791_));
 NAND2_X1 _25263_ (.A1(_07531_),
    .A2(_07791_),
    .ZN(_07792_));
 OR2_X1 _25264_ (.A1(_07513_),
    .A2(_07787_),
    .ZN(_07793_));
 INV_X1 _25265_ (.A(_05482_),
    .ZN(_07794_));
 OAI21_X1 _25266_ (.A(_07792_),
    .B1(_07793_),
    .B2(_07794_),
    .ZN(_07795_));
 AOI21_X1 _25267_ (.A(_07789_),
    .B1(_07795_),
    .B2(_07779_),
    .ZN(_01717_));
 NAND2_X1 _25268_ (.A1(_05482_),
    .A2(_07784_),
    .ZN(_07796_));
 NAND2_X1 _25269_ (.A1(_07737_),
    .A2(_07796_),
    .ZN(_07797_));
 AOI21_X1 _25270_ (.A(_05536_),
    .B1(_07767_),
    .B2(_07797_),
    .ZN(_07798_));
 MUX2_X1 _25271_ (.A(_15526_),
    .B(_07477_),
    .S(_15872_),
    .Z(_07799_));
 OAI22_X4 _25272_ (.A1(_15868_),
    .A2(_05540_),
    .B1(_07799_),
    .B2(_07481_),
    .ZN(_07800_));
 NAND2_X1 _25273_ (.A1(_07526_),
    .A2(_07800_),
    .ZN(_07801_));
 NAND3_X1 _25274_ (.A1(_05482_),
    .A2(_05536_),
    .A3(_07784_),
    .ZN(_07802_));
 OAI21_X1 _25275_ (.A(_07801_),
    .B1(_07802_),
    .B2(_07590_),
    .ZN(_07803_));
 AOI21_X1 _25276_ (.A(_07798_),
    .B1(_07803_),
    .B2(_07779_),
    .ZN(_01718_));
 NAND4_X2 _25277_ (.A1(_05404_),
    .A2(_05457_),
    .A3(_07776_),
    .A4(_07764_),
    .ZN(_07804_));
 NAND2_X1 _25278_ (.A1(_05482_),
    .A2(_05536_),
    .ZN(_07805_));
 OAI21_X1 _25279_ (.A(_07680_),
    .B1(_07804_),
    .B2(_07805_),
    .ZN(_07806_));
 AOI21_X1 _25280_ (.A(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .B1(_07767_),
    .B2(_07806_),
    .ZN(_07807_));
 MUX2_X1 _25281_ (.A(_07532_),
    .B(_07476_),
    .S(_15881_),
    .Z(_07808_));
 NOR2_X1 _25282_ (.A1(_07534_),
    .A2(_07808_),
    .ZN(_07809_));
 AOI21_X4 _25283_ (.A(_07809_),
    .B1(_05577_),
    .B2(_15881_),
    .ZN(_07810_));
 NAND3_X2 _25284_ (.A1(_05482_),
    .A2(_05536_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .ZN(_07811_));
 OAI22_X1 _25285_ (.A1(_07711_),
    .A2(_07810_),
    .B1(_07811_),
    .B2(_07793_),
    .ZN(_07812_));
 AOI21_X1 _25286_ (.A(_07807_),
    .B1(_07812_),
    .B2(_07779_),
    .ZN(_01719_));
 NAND3_X1 _25287_ (.A1(_05459_),
    .A2(_05494_),
    .A3(_07514_),
    .ZN(_07813_));
 NOR3_X2 _25288_ (.A1(_07538_),
    .A2(_07772_),
    .A3(_07813_),
    .ZN(_07814_));
 NAND2_X1 _25289_ (.A1(_07814_),
    .A2(_07774_),
    .ZN(_07815_));
 NOR3_X1 _25290_ (.A1(_07815_),
    .A2(_07705_),
    .A3(_07741_),
    .ZN(_07816_));
 NAND4_X2 _25291_ (.A1(_05404_),
    .A2(_05457_),
    .A3(_07816_),
    .A4(_07764_),
    .ZN(_07817_));
 OAI21_X1 _25292_ (.A(_07528_),
    .B1(_07817_),
    .B2(_07811_),
    .ZN(_07818_));
 AOI21_X1 _25293_ (.A(_05609_),
    .B1(_07758_),
    .B2(_07818_),
    .ZN(_07819_));
 MUX2_X1 _25294_ (.A(_15526_),
    .B(_07477_),
    .S(_15889_),
    .Z(_07820_));
 OAI22_X4 _25295_ (.A1(_15885_),
    .A2(_05611_),
    .B1(_07820_),
    .B2(_07481_),
    .ZN(_07821_));
 NAND2_X1 _25296_ (.A1(_07531_),
    .A2(_07821_),
    .ZN(_07822_));
 AND3_X1 _25297_ (.A1(_05482_),
    .A2(_05536_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .ZN(_07823_));
 NAND3_X2 _25298_ (.A1(_05609_),
    .A2(_07784_),
    .A3(_07823_),
    .ZN(_07824_));
 OR2_X1 _25299_ (.A1(_07537_),
    .A2(_07824_),
    .ZN(_07825_));
 AOI21_X1 _25300_ (.A(_07762_),
    .B1(_07822_),
    .B2(_07825_),
    .ZN(_07826_));
 NOR2_X1 _25301_ (.A1(_07819_),
    .A2(_07826_),
    .ZN(_01720_));
 MUX2_X1 _25302_ (.A(_07477_),
    .B(_15526_),
    .S(_15893_),
    .Z(_07827_));
 OAI22_X4 _25303_ (.A1(_15893_),
    .A2(_05639_),
    .B1(_07827_),
    .B2(_07481_),
    .ZN(_07828_));
 NAND2_X1 _25304_ (.A1(_07531_),
    .A2(_07828_),
    .ZN(_07829_));
 NAND2_X1 _25305_ (.A1(_05609_),
    .A2(_07823_),
    .ZN(_07830_));
 NOR2_X1 _25306_ (.A1(_07787_),
    .A2(_07830_),
    .ZN(_07831_));
 NAND3_X1 _25307_ (.A1(_05625_),
    .A2(_07550_),
    .A3(_07831_),
    .ZN(_07832_));
 AOI21_X1 _25308_ (.A(_07762_),
    .B1(_07829_),
    .B2(_07832_),
    .ZN(_07833_));
 OAI21_X1 _25309_ (.A(_07758_),
    .B1(_07831_),
    .B2(_07590_),
    .ZN(_07834_));
 INV_X1 _25310_ (.A(_05625_),
    .ZN(_07835_));
 AOI21_X1 _25311_ (.A(_07833_),
    .B1(_07834_),
    .B2(_07835_),
    .ZN(_01721_));
 NAND3_X1 _25312_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_05459_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .ZN(_07836_));
 NAND2_X1 _25313_ (.A1(_07737_),
    .A2(_07836_),
    .ZN(_07837_));
 AOI21_X1 _25314_ (.A(_05494_),
    .B1(_07549_),
    .B2(_07837_),
    .ZN(_07838_));
 OAI21_X1 _25315_ (.A(_07792_),
    .B1(_07539_),
    .B2(_07596_),
    .ZN(_07839_));
 AOI21_X1 _25316_ (.A(_07838_),
    .B1(_07839_),
    .B2(_07560_),
    .ZN(_01722_));
 OAI21_X1 _25317_ (.A(_07680_),
    .B1(_07824_),
    .B2(_07835_),
    .ZN(_07840_));
 AOI21_X1 _25318_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B1(_07767_),
    .B2(_07840_),
    .ZN(_07841_));
 MUX2_X1 _25319_ (.A(_07564_),
    .B(_11356_),
    .S(_15901_),
    .Z(_07842_));
 NOR2_X1 _25320_ (.A1(_07480_),
    .A2(_07842_),
    .ZN(_07843_));
 AOI21_X4 _25321_ (.A(_07843_),
    .B1(_05685_),
    .B2(_15905_),
    .ZN(_07844_));
 OR2_X1 _25322_ (.A1(_07563_),
    .A2(_07844_),
    .ZN(_07845_));
 NAND2_X1 _25323_ (.A1(_05625_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .ZN(_07846_));
 OAI21_X1 _25324_ (.A(_07845_),
    .B1(_07846_),
    .B2(_07825_),
    .ZN(_07847_));
 AOI21_X1 _25325_ (.A(_07841_),
    .B1(_07847_),
    .B2(_07779_),
    .ZN(_01723_));
 OR2_X1 _25326_ (.A1(_07787_),
    .A2(_07830_),
    .ZN(_07848_));
 OAI21_X1 _25327_ (.A(_07680_),
    .B1(_07848_),
    .B2(_07846_),
    .ZN(_07849_));
 AOI21_X1 _25328_ (.A(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .B1(_07767_),
    .B2(_07849_),
    .ZN(_07850_));
 MUX2_X1 _25329_ (.A(_11356_),
    .B(_07564_),
    .S(_15913_),
    .Z(_07851_));
 NOR2_X1 _25330_ (.A1(_07480_),
    .A2(_07851_),
    .ZN(_07852_));
 AOI21_X2 _25331_ (.A(_07852_),
    .B1(_05718_),
    .B2(_15913_),
    .ZN(_07853_));
 BUF_X4 _25332_ (.A(_07853_),
    .Z(_07854_));
 NAND3_X4 _25333_ (.A1(_05625_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .ZN(_07855_));
 NAND2_X1 _25334_ (.A1(_07550_),
    .A2(_07831_),
    .ZN(_07856_));
 OAI22_X1 _25335_ (.A1(_07711_),
    .A2(_07854_),
    .B1(_07855_),
    .B2(_07856_),
    .ZN(_07857_));
 AOI21_X1 _25336_ (.A(_07850_),
    .B1(_07857_),
    .B2(_07779_),
    .ZN(_01724_));
 INV_X1 _25337_ (.A(_05742_),
    .ZN(_07858_));
 INV_X1 _25338_ (.A(_05609_),
    .ZN(_07859_));
 NOR4_X4 _25339_ (.A1(_07859_),
    .A2(_07817_),
    .A3(_07811_),
    .A4(_07855_),
    .ZN(_07860_));
 OAI21_X1 _25340_ (.A(_07767_),
    .B1(_07860_),
    .B2(_07596_),
    .ZN(_07861_));
 NAND2_X1 _25341_ (.A1(_07531_),
    .A2(_07524_),
    .ZN(_07862_));
 NAND2_X1 _25342_ (.A1(_07502_),
    .A2(_07860_),
    .ZN(_07863_));
 OAI21_X1 _25343_ (.A(_07862_),
    .B1(_07863_),
    .B2(_07858_),
    .ZN(_07864_));
 AOI22_X1 _25344_ (.A1(_07858_),
    .A2(_07861_),
    .B1(_07864_),
    .B2(_07758_),
    .ZN(_01725_));
 NOR2_X2 _25345_ (.A1(_07848_),
    .A2(_07855_),
    .ZN(_07865_));
 NAND2_X1 _25346_ (.A1(_05742_),
    .A2(_07865_),
    .ZN(_07866_));
 NAND2_X1 _25347_ (.A1(_07528_),
    .A2(_07866_),
    .ZN(_07867_));
 AOI21_X1 _25348_ (.A(_05786_),
    .B1(_07758_),
    .B2(_07867_),
    .ZN(_07868_));
 NAND4_X1 _25349_ (.A1(_05786_),
    .A2(_05742_),
    .A3(_07636_),
    .A4(_07865_),
    .ZN(_07869_));
 AOI21_X1 _25350_ (.A(_07762_),
    .B1(_07869_),
    .B2(_07536_),
    .ZN(_07870_));
 NOR2_X1 _25351_ (.A1(_07868_),
    .A2(_07870_),
    .ZN(_01726_));
 CLKBUF_X3 _25352_ (.A(_07757_),
    .Z(_07871_));
 NAND3_X1 _25353_ (.A1(_05786_),
    .A2(_05742_),
    .A3(_07860_),
    .ZN(_07872_));
 NAND2_X1 _25354_ (.A1(_07737_),
    .A2(_07872_),
    .ZN(_07873_));
 AOI21_X1 _25355_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B1(_07871_),
    .B2(_07873_),
    .ZN(_07874_));
 AND3_X2 _25356_ (.A1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .A2(_05786_),
    .A3(_05742_),
    .ZN(_07875_));
 INV_X1 _25357_ (.A(_07875_),
    .ZN(_07876_));
 OAI21_X1 _25358_ (.A(_07555_),
    .B1(_07863_),
    .B2(_07876_),
    .ZN(_07877_));
 AOI21_X1 _25359_ (.A(_07874_),
    .B1(_07877_),
    .B2(_07779_),
    .ZN(_01727_));
 NAND2_X1 _25360_ (.A1(_07865_),
    .A2(_07875_),
    .ZN(_07878_));
 NAND2_X1 _25361_ (.A1(_07528_),
    .A2(_07878_),
    .ZN(_07879_));
 AOI21_X1 _25362_ (.A(_05875_),
    .B1(_07758_),
    .B2(_07879_),
    .ZN(_07880_));
 NAND4_X1 _25363_ (.A1(_05875_),
    .A2(_07636_),
    .A3(_07865_),
    .A4(_07875_),
    .ZN(_07881_));
 AOI21_X1 _25364_ (.A(_07762_),
    .B1(_07881_),
    .B2(_07570_),
    .ZN(_07882_));
 NOR2_X1 _25365_ (.A1(_07880_),
    .A2(_07882_),
    .ZN(_01728_));
 NAND3_X1 _25366_ (.A1(_05875_),
    .A2(_07860_),
    .A3(_07875_),
    .ZN(_07883_));
 NAND2_X1 _25367_ (.A1(_07737_),
    .A2(_07883_),
    .ZN(_07884_));
 AOI21_X1 _25368_ (.A(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .B1(_07871_),
    .B2(_07884_),
    .ZN(_07885_));
 NAND3_X4 _25369_ (.A1(_05875_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A3(_07875_),
    .ZN(_07886_));
 OAI21_X1 _25370_ (.A(_07580_),
    .B1(_07863_),
    .B2(_07886_),
    .ZN(_07887_));
 AOI21_X1 _25371_ (.A(_07885_),
    .B1(_07887_),
    .B2(_07779_),
    .ZN(_01729_));
 NOR3_X2 _25372_ (.A1(_07848_),
    .A2(_07855_),
    .A3(_07886_),
    .ZN(_07888_));
 NAND3_X1 _25373_ (.A1(_05966_),
    .A2(_07636_),
    .A3(_07888_),
    .ZN(_07889_));
 AOI21_X1 _25374_ (.A(_07762_),
    .B1(_07889_),
    .B2(_07586_),
    .ZN(_07890_));
 NOR4_X2 _25375_ (.A1(_07804_),
    .A2(_07830_),
    .A3(_07855_),
    .A4(_07886_),
    .ZN(_07891_));
 OAI21_X1 _25376_ (.A(_07767_),
    .B1(_07891_),
    .B2(_07596_),
    .ZN(_07892_));
 INV_X1 _25377_ (.A(_05966_),
    .ZN(_07893_));
 AOI21_X1 _25378_ (.A(_07890_),
    .B1(_07892_),
    .B2(_07893_),
    .ZN(_01730_));
 AND3_X1 _25379_ (.A1(_05875_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A3(_07875_),
    .ZN(_07894_));
 NAND3_X1 _25380_ (.A1(_05966_),
    .A2(_07860_),
    .A3(_07894_),
    .ZN(_07895_));
 NAND2_X1 _25381_ (.A1(_07737_),
    .A2(_07895_),
    .ZN(_07896_));
 AOI21_X1 _25382_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .B1(_07871_),
    .B2(_07896_),
    .ZN(_07897_));
 NAND4_X1 _25383_ (.A1(_05966_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .A3(_07860_),
    .A4(_07894_),
    .ZN(_07898_));
 OAI21_X1 _25384_ (.A(_07601_),
    .B1(_07898_),
    .B2(_07596_),
    .ZN(_07899_));
 AOI21_X1 _25385_ (.A(_07897_),
    .B1(_07899_),
    .B2(_07779_),
    .ZN(_01731_));
 AND2_X2 _25386_ (.A1(_05966_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .ZN(_07900_));
 NAND2_X1 _25387_ (.A1(_07888_),
    .A2(_07900_),
    .ZN(_07901_));
 NAND2_X1 _25388_ (.A1(_07737_),
    .A2(_07901_),
    .ZN(_07902_));
 AOI21_X1 _25389_ (.A(_06034_),
    .B1(_07871_),
    .B2(_07902_),
    .ZN(_07903_));
 NAND4_X1 _25390_ (.A1(_06034_),
    .A2(_07502_),
    .A3(_07888_),
    .A4(_07900_),
    .ZN(_07904_));
 NAND2_X1 _25391_ (.A1(_07606_),
    .A2(_07904_),
    .ZN(_07905_));
 AOI21_X1 _25392_ (.A(_07903_),
    .B1(_07905_),
    .B2(_07779_),
    .ZN(_01732_));
 NAND2_X1 _25393_ (.A1(_07528_),
    .A2(_07813_),
    .ZN(_07906_));
 AOI21_X1 _25394_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B1(_07560_),
    .B2(_07906_),
    .ZN(_07907_));
 NAND3_X1 _25395_ (.A1(_07514_),
    .A2(_07504_),
    .A3(_07515_),
    .ZN(_07908_));
 AOI21_X1 _25396_ (.A(_07509_),
    .B1(_07801_),
    .B2(_07908_),
    .ZN(_07909_));
 NOR2_X1 _25397_ (.A1(_07907_),
    .A2(_07909_),
    .ZN(_01733_));
 INV_X1 _25398_ (.A(_06091_),
    .ZN(_07910_));
 NAND2_X1 _25399_ (.A1(_06034_),
    .A2(_07900_),
    .ZN(_07911_));
 NOR4_X4 _25400_ (.A1(_07824_),
    .A2(_07855_),
    .A3(_07886_),
    .A4(_07911_),
    .ZN(_07912_));
 OAI21_X1 _25401_ (.A(_07767_),
    .B1(_07912_),
    .B2(_07596_),
    .ZN(_07913_));
 INV_X2 _25402_ (.A(_07616_),
    .ZN(_07914_));
 NAND2_X1 _25403_ (.A1(_07502_),
    .A2(_07912_),
    .ZN(_07915_));
 OAI22_X1 _25404_ (.A1(_07711_),
    .A2(_07914_),
    .B1(_07915_),
    .B2(_07910_),
    .ZN(_07916_));
 AOI22_X1 _25405_ (.A1(_07910_),
    .A2(_07913_),
    .B1(_07916_),
    .B2(_07758_),
    .ZN(_01734_));
 NAND3_X1 _25406_ (.A1(_06034_),
    .A2(_07891_),
    .A3(_07900_),
    .ZN(_07917_));
 OAI21_X1 _25407_ (.A(_07680_),
    .B1(_07917_),
    .B2(_07910_),
    .ZN(_07918_));
 AOI21_X1 _25408_ (.A(_06120_),
    .B1(_07871_),
    .B2(_07918_),
    .ZN(_07919_));
 NAND2_X1 _25409_ (.A1(_06091_),
    .A2(_06120_),
    .ZN(_07920_));
 OAI21_X1 _25410_ (.A(_07625_),
    .B1(_07904_),
    .B2(_07920_),
    .ZN(_07921_));
 CLKBUF_X3 _25411_ (.A(_07757_),
    .Z(_07922_));
 AOI21_X1 _25412_ (.A(_07919_),
    .B1(_07921_),
    .B2(_07922_),
    .ZN(_01735_));
 NAND4_X2 _25413_ (.A1(_06034_),
    .A2(_07860_),
    .A3(_07894_),
    .A4(_07900_),
    .ZN(_07923_));
 OAI21_X1 _25414_ (.A(_07680_),
    .B1(_07923_),
    .B2(_07920_),
    .ZN(_07924_));
 AOI21_X1 _25415_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B1(_07871_),
    .B2(_07924_),
    .ZN(_07925_));
 NAND3_X2 _25416_ (.A1(_06091_),
    .A2(_06120_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .ZN(_07926_));
 OAI21_X1 _25417_ (.A(_07641_),
    .B1(_07915_),
    .B2(_07926_),
    .ZN(_07927_));
 AOI21_X1 _25418_ (.A(_07925_),
    .B1(_07927_),
    .B2(_07922_),
    .ZN(_01736_));
 INV_X1 _25419_ (.A(_06034_),
    .ZN(_07928_));
 NOR3_X2 _25420_ (.A1(_07928_),
    .A2(_07901_),
    .A3(_07926_),
    .ZN(_07929_));
 NAND3_X1 _25421_ (.A1(_06193_),
    .A2(_07636_),
    .A3(_07929_),
    .ZN(_07930_));
 AOI21_X1 _25422_ (.A(_07762_),
    .B1(_07930_),
    .B2(_07652_),
    .ZN(_07931_));
 AND3_X1 _25423_ (.A1(_06091_),
    .A2(_06120_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .ZN(_07932_));
 NAND4_X1 _25424_ (.A1(_06034_),
    .A2(_07891_),
    .A3(_07900_),
    .A4(_07932_),
    .ZN(_07933_));
 NAND2_X1 _25425_ (.A1(_07711_),
    .A2(_07933_),
    .ZN(_07934_));
 NAND2_X1 _25426_ (.A1(_07758_),
    .A2(_07934_),
    .ZN(_07935_));
 INV_X1 _25427_ (.A(_06193_),
    .ZN(_07936_));
 AOI21_X1 _25428_ (.A(_07931_),
    .B1(_07935_),
    .B2(_07936_),
    .ZN(_01737_));
 NOR3_X2 _25429_ (.A1(_07936_),
    .A2(_07923_),
    .A3(_07926_),
    .ZN(_07937_));
 NAND3_X2 _25430_ (.A1(_04547_),
    .A2(_07563_),
    .A3(_07937_),
    .ZN(_07938_));
 AOI21_X1 _25431_ (.A(_07762_),
    .B1(_07938_),
    .B2(_07658_),
    .ZN(_07939_));
 OAI21_X1 _25432_ (.A(_07767_),
    .B1(_07937_),
    .B2(_07596_),
    .ZN(_07940_));
 INV_X1 _25433_ (.A(_04547_),
    .ZN(_07941_));
 AOI21_X1 _25434_ (.A(_07939_),
    .B1(_07940_),
    .B2(_07941_),
    .ZN(_01738_));
 OR3_X2 _25435_ (.A1(_07936_),
    .A2(_07941_),
    .A3(_07933_),
    .ZN(_07942_));
 NAND2_X1 _25436_ (.A1(_07737_),
    .A2(_07942_),
    .ZN(_07943_));
 AOI21_X1 _25437_ (.A(_04751_),
    .B1(_07871_),
    .B2(_07943_),
    .ZN(_07944_));
 NAND4_X2 _25438_ (.A1(_06193_),
    .A2(_04547_),
    .A3(_07563_),
    .A4(_07929_),
    .ZN(_07945_));
 INV_X1 _25439_ (.A(_04751_),
    .ZN(_07946_));
 OAI21_X1 _25440_ (.A(_07670_),
    .B1(_07945_),
    .B2(_07946_),
    .ZN(_07947_));
 AOI21_X1 _25441_ (.A(_07944_),
    .B1(_07947_),
    .B2(_07922_),
    .ZN(_01739_));
 NAND4_X2 _25442_ (.A1(_06193_),
    .A2(_04547_),
    .A3(_07912_),
    .A4(_07932_),
    .ZN(_07948_));
 OAI21_X1 _25443_ (.A(_07680_),
    .B1(_07948_),
    .B2(_07946_),
    .ZN(_07949_));
 AOI21_X1 _25444_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B1(_07871_),
    .B2(_07949_),
    .ZN(_07950_));
 NAND2_X1 _25445_ (.A1(_04751_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .ZN(_07951_));
 OAI21_X1 _25446_ (.A(_07677_),
    .B1(_07938_),
    .B2(_07951_),
    .ZN(_07952_));
 AOI21_X1 _25447_ (.A(_07950_),
    .B1(_07952_),
    .B2(_07922_),
    .ZN(_01740_));
 OAI21_X1 _25448_ (.A(_07680_),
    .B1(_07942_),
    .B2(_07951_),
    .ZN(_07953_));
 AOI21_X1 _25449_ (.A(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .B1(_07871_),
    .B2(_07953_),
    .ZN(_07954_));
 NAND3_X2 _25450_ (.A1(_04751_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .ZN(_07955_));
 OAI21_X1 _25451_ (.A(_07690_),
    .B1(_07945_),
    .B2(_07955_),
    .ZN(_07956_));
 AOI21_X1 _25452_ (.A(_07954_),
    .B1(_07956_),
    .B2(_07922_),
    .ZN(_01741_));
 OAI21_X1 _25453_ (.A(_07680_),
    .B1(_07948_),
    .B2(_07955_),
    .ZN(_07957_));
 AOI21_X1 _25454_ (.A(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .B1(_07871_),
    .B2(_07957_),
    .ZN(_07958_));
 INV_X1 _25455_ (.A(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .ZN(_07959_));
 OR2_X1 _25456_ (.A1(_07959_),
    .A2(_07955_),
    .ZN(_07960_));
 OAI21_X1 _25457_ (.A(_07697_),
    .B1(_07938_),
    .B2(_07960_),
    .ZN(_07961_));
 AOI21_X1 _25458_ (.A(_07958_),
    .B1(_07961_),
    .B2(_07922_),
    .ZN(_01742_));
 OAI21_X1 _25459_ (.A(_07680_),
    .B1(_07942_),
    .B2(_07960_),
    .ZN(_07962_));
 AOI21_X1 _25460_ (.A(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .B1(_07757_),
    .B2(_07962_),
    .ZN(_07963_));
 NAND2_X1 _25461_ (.A1(_07526_),
    .A2(_07709_),
    .ZN(_07964_));
 NOR2_X1 _25462_ (.A1(_07959_),
    .A2(_07955_),
    .ZN(_07965_));
 NAND2_X1 _25463_ (.A1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .A2(_07965_),
    .ZN(_07966_));
 OAI21_X1 _25464_ (.A(_07964_),
    .B1(_07945_),
    .B2(_07966_),
    .ZN(_07967_));
 AOI21_X1 _25465_ (.A(_07963_),
    .B1(_07967_),
    .B2(_07922_),
    .ZN(_01743_));
 NAND2_X1 _25466_ (.A1(_07504_),
    .A2(_07773_),
    .ZN(_07968_));
 OAI21_X1 _25467_ (.A(_07968_),
    .B1(_07810_),
    .B2(_07711_),
    .ZN(_07969_));
 OAI21_X1 _25468_ (.A(_07507_),
    .B1(_07540_),
    .B2(_07596_),
    .ZN(_07970_));
 AOI22_X1 _25469_ (.A1(_07559_),
    .A2(_07969_),
    .B1(_07970_),
    .B2(_07772_),
    .ZN(_01744_));
 OAI21_X1 _25470_ (.A(_07502_),
    .B1(_07948_),
    .B2(_07966_),
    .ZN(_07971_));
 AOI21_X1 _25471_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B1(_07757_),
    .B2(_07971_),
    .ZN(_07972_));
 AND2_X1 _25472_ (.A1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .A2(_07965_),
    .ZN(_07973_));
 NAND2_X1 _25473_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_07973_),
    .ZN(_07974_));
 OAI21_X1 _25474_ (.A(_07719_),
    .B1(_07938_),
    .B2(_07974_),
    .ZN(_07975_));
 AOI21_X1 _25475_ (.A(_07972_),
    .B1(_07975_),
    .B2(_07922_),
    .ZN(_01745_));
 OAI21_X1 _25476_ (.A(_07502_),
    .B1(_07942_),
    .B2(_07974_),
    .ZN(_07976_));
 AOI21_X1 _25477_ (.A(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .B1(_07757_),
    .B2(_07976_),
    .ZN(_07977_));
 AND2_X1 _25478_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_07973_),
    .ZN(_07978_));
 NAND2_X1 _25479_ (.A1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A2(_07978_),
    .ZN(_07979_));
 OAI21_X1 _25480_ (.A(_07729_),
    .B1(_07945_),
    .B2(_07979_),
    .ZN(_07980_));
 AOI21_X1 _25481_ (.A(_07977_),
    .B1(_07980_),
    .B2(_07922_),
    .ZN(_01746_));
 OAI21_X1 _25482_ (.A(_07502_),
    .B1(_07948_),
    .B2(_07979_),
    .ZN(_07981_));
 AOI21_X1 _25483_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B1(_07757_),
    .B2(_07981_),
    .ZN(_07982_));
 BUF_X4 _25484_ (.A(_07745_),
    .Z(_07983_));
 NAND2_X1 _25485_ (.A1(_07526_),
    .A2(_07983_),
    .ZN(_07984_));
 NAND3_X1 _25486_ (.A1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .A3(_07978_),
    .ZN(_07985_));
 OAI21_X1 _25487_ (.A(_07984_),
    .B1(_07938_),
    .B2(_07985_),
    .ZN(_07986_));
 AOI21_X1 _25488_ (.A(_07982_),
    .B1(_07986_),
    .B2(_07922_),
    .ZN(_01747_));
 OAI21_X1 _25489_ (.A(_07502_),
    .B1(_07942_),
    .B2(_07985_),
    .ZN(_07987_));
 AOI21_X1 _25490_ (.A(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .B1(_07757_),
    .B2(_07987_),
    .ZN(_07988_));
 NOR2_X1 _25491_ (.A1(_07942_),
    .A2(_07985_),
    .ZN(_07989_));
 NAND3_X1 _25492_ (.A1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .A2(_07528_),
    .A3(_07989_),
    .ZN(_07990_));
 NAND2_X1 _25493_ (.A1(_07749_),
    .A2(_07990_),
    .ZN(_07991_));
 AOI21_X1 _25494_ (.A(_07988_),
    .B1(_07991_),
    .B2(_07758_),
    .ZN(_01748_));
 NAND2_X1 _25495_ (.A1(_07636_),
    .A2(_07814_),
    .ZN(_07992_));
 INV_X1 _25496_ (.A(_05606_),
    .ZN(_07993_));
 OAI21_X1 _25497_ (.A(_07822_),
    .B1(_07992_),
    .B2(_07993_),
    .ZN(_07994_));
 OAI21_X1 _25498_ (.A(_07507_),
    .B1(_07814_),
    .B2(_07526_),
    .ZN(_07995_));
 AOI22_X1 _25499_ (.A1(_07559_),
    .A2(_07994_),
    .B1(_07995_),
    .B2(_07993_),
    .ZN(_01749_));
 NAND4_X1 _25500_ (.A1(_05606_),
    .A2(_05628_),
    .A3(_07636_),
    .A4(_07773_),
    .ZN(_07996_));
 AOI21_X1 _25501_ (.A(_07509_),
    .B1(_07829_),
    .B2(_07996_),
    .ZN(_07997_));
 OAI21_X1 _25502_ (.A(_07504_),
    .B1(_07541_),
    .B2(_07993_),
    .ZN(_07998_));
 AOI21_X1 _25503_ (.A(_05628_),
    .B1(_07546_),
    .B2(_07998_),
    .ZN(_07999_));
 NOR2_X1 _25504_ (.A1(_07997_),
    .A2(_07999_),
    .ZN(_01750_));
 NAND3_X1 _25505_ (.A1(_05606_),
    .A2(_05628_),
    .A3(_07814_),
    .ZN(_08000_));
 NAND2_X1 _25506_ (.A1(_07636_),
    .A2(_08000_),
    .ZN(_08001_));
 AOI21_X1 _25507_ (.A(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .B1(_07507_),
    .B2(_08001_),
    .ZN(_08002_));
 OAI21_X1 _25508_ (.A(_07845_),
    .B1(_07992_),
    .B2(_07518_),
    .ZN(_08003_));
 AOI21_X1 _25509_ (.A(_08002_),
    .B1(_08003_),
    .B2(_07560_),
    .ZN(_01751_));
 OR2_X1 _25510_ (.A1(_07518_),
    .A2(_07541_),
    .ZN(_08004_));
 NAND2_X1 _25511_ (.A1(_07636_),
    .A2(_08004_),
    .ZN(_08005_));
 AOI21_X1 _25512_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .B1(_07507_),
    .B2(_08005_),
    .ZN(_08006_));
 OR3_X1 _25513_ (.A1(_07517_),
    .A2(_07513_),
    .A3(_08004_),
    .ZN(_08007_));
 OAI21_X1 _25514_ (.A(_08007_),
    .B1(_07854_),
    .B2(_07711_),
    .ZN(_08008_));
 AOI21_X1 _25515_ (.A(_08006_),
    .B1(_08008_),
    .B2(_07560_),
    .ZN(_01752_));
 NOR4_X1 _25516_ (.A1(_05241_),
    .A2(_05292_),
    .A3(_05303_),
    .A4(_05286_),
    .ZN(_08009_));
 NOR3_X1 _25517_ (.A1(_05241_),
    .A2(_05292_),
    .A3(_05286_),
    .ZN(_08010_));
 NAND2_X1 _25518_ (.A1(_03398_),
    .A2(_03399_),
    .ZN(_08011_));
 AOI21_X1 _25519_ (.A(_08009_),
    .B1(_08010_),
    .B2(_08011_),
    .ZN(_08012_));
 NAND2_X1 _25520_ (.A1(_05241_),
    .A2(_05304_),
    .ZN(_08013_));
 OAI221_X1 _25521_ (.A(_08012_),
    .B1(_08013_),
    .B2(_05311_),
    .C1(_05286_),
    .C2(_05282_),
    .ZN(_08014_));
 AND3_X1 _25522_ (.A1(_05241_),
    .A2(_05311_),
    .A3(_05297_),
    .ZN(_08015_));
 NAND2_X1 _25523_ (.A1(_05283_),
    .A2(_05297_),
    .ZN(_08016_));
 NOR3_X1 _25524_ (.A1(_05292_),
    .A2(_08011_),
    .A3(_08016_),
    .ZN(_08017_));
 NOR3_X1 _25525_ (.A1(net274),
    .A2(_05289_),
    .A3(_08016_),
    .ZN(_08018_));
 OR3_X1 _25526_ (.A1(_08015_),
    .A2(_08017_),
    .A3(_08018_),
    .ZN(_08019_));
 NAND2_X1 _25527_ (.A1(_10895_),
    .A2(_05316_),
    .ZN(_08020_));
 NOR4_X1 _25528_ (.A1(_03645_),
    .A2(_08014_),
    .A3(_08019_),
    .A4(_08020_),
    .ZN(_08021_));
 MUX2_X1 _25529_ (.A(_05315_),
    .B(_08021_),
    .S(_06248_),
    .Z(_08022_));
 OAI22_X2 _25530_ (.A1(net308),
    .A2(_05314_),
    .B1(_05316_),
    .B2(_06249_),
    .ZN(_08023_));
 OAI21_X2 _25531_ (.A(_03886_),
    .B1(_08022_),
    .B2(_08023_),
    .ZN(_08024_));
 XNOR2_X1 _25532_ (.A(_15846_),
    .B(_15860_),
    .ZN(_08025_));
 NOR2_X1 _25533_ (.A1(_11066_),
    .A2(_15853_),
    .ZN(_08026_));
 AOI22_X1 _25534_ (.A1(_11066_),
    .A2(_03594_),
    .B1(_08025_),
    .B2(_08026_),
    .ZN(_08027_));
 OR4_X2 _25535_ (.A1(_15509_),
    .A2(_15513_),
    .A3(_15841_),
    .A4(_08027_),
    .ZN(_08028_));
 OR3_X2 _25536_ (.A1(_07617_),
    .A2(_07619_),
    .A3(_08028_),
    .ZN(_08029_));
 NAND2_X1 _25537_ (.A1(_03435_),
    .A2(_01159_),
    .ZN(_08030_));
 NOR3_X2 _25538_ (.A1(_10742_),
    .A2(_03471_),
    .A3(_03608_),
    .ZN(_08031_));
 NOR4_X4 _25539_ (.A1(_06262_),
    .A2(_06272_),
    .A3(_08030_),
    .A4(_08031_),
    .ZN(_08032_));
 AOI21_X1 _25540_ (.A(_07484_),
    .B1(_03485_),
    .B2(_03487_),
    .ZN(_08033_));
 OAI21_X1 _25541_ (.A(_08033_),
    .B1(_03603_),
    .B2(_04608_),
    .ZN(_08034_));
 NAND2_X1 _25542_ (.A1(_03518_),
    .A2(_08034_),
    .ZN(_08035_));
 AND3_X1 _25543_ (.A1(_03439_),
    .A2(_08032_),
    .A3(_08035_),
    .ZN(_08036_));
 AND3_X1 _25544_ (.A1(_08024_),
    .A2(_08029_),
    .A3(_08036_),
    .ZN(_08037_));
 CLKBUF_X3 _25545_ (.A(_08037_),
    .Z(_08038_));
 INV_X1 _25546_ (.A(_08029_),
    .ZN(_08039_));
 AND2_X1 _25547_ (.A1(_04756_),
    .A2(_08039_),
    .ZN(_08040_));
 BUF_X2 _25548_ (.A(_08040_),
    .Z(_08041_));
 OR3_X1 _25549_ (.A1(\cs_registers_i.mhpmcounter[2][0] ),
    .A2(_08038_),
    .A3(_08041_),
    .ZN(_08042_));
 OR2_X2 _25550_ (.A1(_07487_),
    .A2(_08028_),
    .ZN(_08043_));
 OR2_X2 _25551_ (.A1(_07511_),
    .A2(_08043_),
    .ZN(_08044_));
 NOR2_X4 _25552_ (.A1(_05745_),
    .A2(_08044_),
    .ZN(_08045_));
 CLKBUF_X3 _25553_ (.A(_08045_),
    .Z(_08046_));
 CLKBUF_X3 _25554_ (.A(_08046_),
    .Z(_08047_));
 NOR2_X4 _25555_ (.A1(_07511_),
    .A2(_08043_),
    .ZN(_08048_));
 AOI211_X2 _25556_ (.A(net307),
    .B(_06251_),
    .C1(_05314_),
    .C2(_05338_),
    .ZN(_08049_));
 NAND3_X4 _25557_ (.A1(_03439_),
    .A2(_04261_),
    .A3(_08032_),
    .ZN(_08050_));
 NOR3_X2 _25558_ (.A1(_08048_),
    .A2(net378),
    .A3(_08050_),
    .ZN(_08051_));
 CLKBUF_X3 _25559_ (.A(_08051_),
    .Z(_08052_));
 AOI22_X1 _25560_ (.A1(_07482_),
    .A2(_08047_),
    .B1(_08052_),
    .B2(_05356_),
    .ZN(_08053_));
 AND2_X1 _25561_ (.A1(_08042_),
    .A2(_08053_),
    .ZN(_01753_));
 NAND2_X2 _25562_ (.A1(_04558_),
    .A2(_08048_),
    .ZN(_08054_));
 CLKBUF_X3 _25563_ (.A(_08054_),
    .Z(_08055_));
 NOR2_X1 _25564_ (.A1(_07525_),
    .A2(_08055_),
    .ZN(_08056_));
 NAND2_X1 _25565_ (.A1(_05750_),
    .A2(_08054_),
    .ZN(_08057_));
 AND4_X1 _25566_ (.A1(_05607_),
    .A2(\cs_registers_i.mhpmcounter[2][7] ),
    .A3(\cs_registers_i.mhpmcounter[2][8] ),
    .A4(\cs_registers_i.mhpmcounter[2][9] ),
    .ZN(_08058_));
 AND3_X1 _25567_ (.A1(\cs_registers_i.mhpmcounter[2][2] ),
    .A2(_15532_),
    .A3(\cs_registers_i.mhpmcounter[2][3] ),
    .ZN(_08059_));
 BUF_X2 _25568_ (.A(_08059_),
    .Z(_08060_));
 AND2_X1 _25569_ (.A1(_05538_),
    .A2(\cs_registers_i.mhpmcounter[2][5] ),
    .ZN(_08061_));
 AND2_X1 _25570_ (.A1(_08060_),
    .A2(_08061_),
    .ZN(_08062_));
 AND2_X1 _25571_ (.A1(_08058_),
    .A2(_08062_),
    .ZN(_08063_));
 AOI21_X1 _25572_ (.A(_08057_),
    .B1(_08063_),
    .B2(_08038_),
    .ZN(_08064_));
 INV_X1 _25573_ (.A(_05750_),
    .ZN(_08065_));
 AND2_X1 _25574_ (.A1(_08058_),
    .A2(_08061_),
    .ZN(_08066_));
 AND4_X1 _25575_ (.A1(_08065_),
    .A2(_08052_),
    .A3(_08060_),
    .A4(_08066_),
    .ZN(_08067_));
 OR3_X1 _25576_ (.A1(_08056_),
    .A2(_08064_),
    .A3(_08067_),
    .ZN(_01754_));
 NOR2_X1 _25577_ (.A1(_05789_),
    .A2(_08046_),
    .ZN(_08068_));
 AND3_X1 _25578_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(\cs_registers_i.mhpmcounter[2][2] ),
    .A3(\cs_registers_i.mhpmcounter[2][0] ),
    .ZN(_08069_));
 AND2_X1 _25579_ (.A1(\cs_registers_i.mhpmcounter[2][3] ),
    .A2(_08069_),
    .ZN(_08070_));
 AND4_X1 _25580_ (.A1(_05750_),
    .A2(_08058_),
    .A3(_08061_),
    .A4(_08070_),
    .ZN(_08071_));
 NAND4_X1 _25581_ (.A1(_08024_),
    .A2(_08029_),
    .A3(_08036_),
    .A4(_08071_),
    .ZN(_08072_));
 MUX2_X1 _25582_ (.A(_05789_),
    .B(_08068_),
    .S(_08072_),
    .Z(_08073_));
 AOI21_X1 _25583_ (.A(_08073_),
    .B1(_08047_),
    .B2(_07535_),
    .ZN(_01755_));
 OR2_X1 _25584_ (.A1(\cs_registers_i.mhpmcounter[2][12] ),
    .A2(_08046_),
    .ZN(_08074_));
 AND4_X1 _25585_ (.A1(_05789_),
    .A2(_05750_),
    .A3(_08058_),
    .A4(_08062_),
    .ZN(_08075_));
 AOI21_X1 _25586_ (.A(_08074_),
    .B1(_08075_),
    .B2(_08037_),
    .ZN(_08076_));
 AND4_X1 _25587_ (.A1(\cs_registers_i.mhpmcounter[2][12] ),
    .A2(_05789_),
    .A3(_05750_),
    .A4(_08066_),
    .ZN(_08077_));
 AND2_X1 _25588_ (.A1(_08060_),
    .A2(_08077_),
    .ZN(_08078_));
 AOI221_X1 _25589_ (.A(_08076_),
    .B1(_08078_),
    .B2(_08038_),
    .C1(_08041_),
    .C2(_07554_),
    .ZN(_01756_));
 NOR2_X1 _25590_ (.A1(_07569_),
    .A2(_08054_),
    .ZN(_08079_));
 BUF_X2 _25591_ (.A(_08070_),
    .Z(_08080_));
 AND4_X1 _25592_ (.A1(_05878_),
    .A2(_08051_),
    .A3(_08080_),
    .A4(_08077_),
    .ZN(_08081_));
 NAND3_X1 _25593_ (.A1(_08052_),
    .A2(_08080_),
    .A3(_08077_),
    .ZN(_08082_));
 CLKBUF_X3 _25594_ (.A(_08046_),
    .Z(_08083_));
 NOR2_X1 _25595_ (.A1(_05878_),
    .A2(_08083_),
    .ZN(_08084_));
 AOI211_X2 _25596_ (.A(_08079_),
    .B(_08081_),
    .C1(_08082_),
    .C2(_08084_),
    .ZN(_01757_));
 OR2_X1 _25597_ (.A1(\cs_registers_i.mhpmcounter[2][14] ),
    .A2(_08046_),
    .ZN(_08085_));
 NAND2_X1 _25598_ (.A1(_08060_),
    .A2(_08077_),
    .ZN(_08086_));
 NOR4_X2 _25599_ (.A1(_08048_),
    .A2(net378),
    .A3(_08050_),
    .A4(_08086_),
    .ZN(_08087_));
 AOI21_X1 _25600_ (.A(_08085_),
    .B1(_08087_),
    .B2(_05878_),
    .ZN(_08088_));
 INV_X1 _25601_ (.A(_07579_),
    .ZN(_08089_));
 AND2_X1 _25602_ (.A1(_05878_),
    .A2(_08087_),
    .ZN(_08090_));
 AOI221_X1 _25603_ (.A(_08088_),
    .B1(_08047_),
    .B2(_08089_),
    .C1(\cs_registers_i.mhpmcounter[2][14] ),
    .C2(_08090_),
    .ZN(_01758_));
 OR2_X1 _25604_ (.A1(\cs_registers_i.mhpmcounter[2][15] ),
    .A2(_08046_),
    .ZN(_08091_));
 AND2_X1 _25605_ (.A1(_05878_),
    .A2(\cs_registers_i.mhpmcounter[2][14] ),
    .ZN(_08092_));
 AND3_X1 _25606_ (.A1(_08080_),
    .A2(_08077_),
    .A3(_08092_),
    .ZN(_08093_));
 AOI21_X1 _25607_ (.A(_08091_),
    .B1(_08093_),
    .B2(_08037_),
    .ZN(_08094_));
 AND4_X1 _25608_ (.A1(\cs_registers_i.mhpmcounter[2][15] ),
    .A2(_08080_),
    .A3(_08077_),
    .A4(_08092_),
    .ZN(_08095_));
 AOI221_X1 _25609_ (.A(_08094_),
    .B1(_08095_),
    .B2(_08038_),
    .C1(_08041_),
    .C2(_07585_),
    .ZN(_01759_));
 OR2_X1 _25610_ (.A1(\cs_registers_i.mhpmcounter[2][16] ),
    .A2(_08045_),
    .ZN(_08096_));
 AND2_X1 _25611_ (.A1(\cs_registers_i.mhpmcounter[2][15] ),
    .A2(_08092_),
    .ZN(_08097_));
 AOI21_X1 _25612_ (.A(_08096_),
    .B1(_08097_),
    .B2(_08087_),
    .ZN(_08098_));
 AND3_X1 _25613_ (.A1(\cs_registers_i.mhpmcounter[2][16] ),
    .A2(_08078_),
    .A3(_08097_),
    .ZN(_08099_));
 INV_X1 _25614_ (.A(_07600_),
    .ZN(_08100_));
 AOI221_X1 _25615_ (.A(_08098_),
    .B1(_08099_),
    .B2(_08038_),
    .C1(_08041_),
    .C2(_08100_),
    .ZN(_01760_));
 AND4_X1 _25616_ (.A1(\cs_registers_i.mhpmcounter[2][16] ),
    .A2(_08070_),
    .A3(_08077_),
    .A4(_08097_),
    .ZN(_08101_));
 INV_X1 _25617_ (.A(_08101_),
    .ZN(_08102_));
 NOR4_X4 _25618_ (.A1(_08048_),
    .A2(net379),
    .A3(_08050_),
    .A4(_08102_),
    .ZN(_08103_));
 NOR3_X1 _25619_ (.A1(_06038_),
    .A2(_08046_),
    .A3(_08103_),
    .ZN(_08104_));
 BUF_X4 _25620_ (.A(_08103_),
    .Z(_08105_));
 AOI221_X1 _25621_ (.A(_08104_),
    .B1(_08083_),
    .B2(_07605_),
    .C1(_06038_),
    .C2(_08105_),
    .ZN(_01761_));
 NAND2_X1 _25622_ (.A1(_06095_),
    .A2(_08055_),
    .ZN(_08106_));
 NAND3_X4 _25623_ (.A1(\cs_registers_i.mhpmcounter[2][16] ),
    .A2(_08078_),
    .A3(_08097_),
    .ZN(_08107_));
 NOR4_X4 _25624_ (.A1(_08048_),
    .A2(net379),
    .A3(_08050_),
    .A4(_08107_),
    .ZN(_08108_));
 AND2_X1 _25625_ (.A1(_06038_),
    .A2(_08108_),
    .ZN(_08109_));
 INV_X1 _25626_ (.A(_06038_),
    .ZN(_08110_));
 NOR4_X1 _25627_ (.A1(_08110_),
    .A2(_06095_),
    .A3(_08048_),
    .A4(_08107_),
    .ZN(_08111_));
 CLKBUF_X3 _25628_ (.A(_08048_),
    .Z(_08112_));
 AOI21_X1 _25629_ (.A(_08111_),
    .B1(_08112_),
    .B2(_07914_),
    .ZN(_08113_));
 NOR2_X2 _25630_ (.A1(_08083_),
    .A2(_08052_),
    .ZN(_08114_));
 OAI22_X1 _25631_ (.A1(_08106_),
    .A2(_08109_),
    .B1(_08113_),
    .B2(_08114_),
    .ZN(_01762_));
 AND2_X1 _25632_ (.A1(_07624_),
    .A2(_08047_),
    .ZN(_08115_));
 OR2_X1 _25633_ (.A1(_06124_),
    .A2(_08046_),
    .ZN(_08116_));
 AND2_X1 _25634_ (.A1(_06038_),
    .A2(_06095_),
    .ZN(_08117_));
 AOI21_X1 _25635_ (.A(_08116_),
    .B1(_08117_),
    .B2(_08105_),
    .ZN(_08118_));
 AND3_X1 _25636_ (.A1(_06124_),
    .A2(_08105_),
    .A3(_08117_),
    .ZN(_08119_));
 NOR3_X1 _25637_ (.A1(_08115_),
    .A2(_08118_),
    .A3(_08119_),
    .ZN(_01763_));
 OR3_X1 _25638_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(_08038_),
    .A3(_08041_),
    .ZN(_08120_));
 INV_X1 _25639_ (.A(_15533_),
    .ZN(_08121_));
 AOI22_X1 _25640_ (.A1(_07635_),
    .A2(_08047_),
    .B1(_08052_),
    .B2(_08121_),
    .ZN(_08122_));
 AND2_X1 _25641_ (.A1(_08120_),
    .A2(_08122_),
    .ZN(_01764_));
 NAND2_X1 _25642_ (.A1(\cs_registers_i.mhpmcounter[2][20] ),
    .A2(_08055_),
    .ZN(_08123_));
 AND3_X1 _25643_ (.A1(_06124_),
    .A2(_08108_),
    .A3(_08117_),
    .ZN(_08124_));
 CLKBUF_X3 _25644_ (.A(_08044_),
    .Z(_08125_));
 NOR2_X1 _25645_ (.A1(_07640_),
    .A2(_08125_),
    .ZN(_08126_));
 NAND2_X1 _25646_ (.A1(_06124_),
    .A2(_08117_),
    .ZN(_08127_));
 NOR3_X1 _25647_ (.A1(\cs_registers_i.mhpmcounter[2][20] ),
    .A2(_08107_),
    .A3(_08127_),
    .ZN(_08128_));
 CLKBUF_X3 _25648_ (.A(_08125_),
    .Z(_08129_));
 AOI21_X1 _25649_ (.A(_08126_),
    .B1(_08128_),
    .B2(_08129_),
    .ZN(_08130_));
 OAI22_X1 _25650_ (.A1(_08123_),
    .A2(_08124_),
    .B1(_08130_),
    .B2(_08114_),
    .ZN(_01765_));
 OR2_X1 _25651_ (.A1(\cs_registers_i.mhpmcounter[2][21] ),
    .A2(_08045_),
    .ZN(_08131_));
 AND4_X1 _25652_ (.A1(_06038_),
    .A2(_06095_),
    .A3(_06124_),
    .A4(\cs_registers_i.mhpmcounter[2][20] ),
    .ZN(_08132_));
 AOI21_X1 _25653_ (.A(_08131_),
    .B1(_08132_),
    .B2(_08105_),
    .ZN(_08133_));
 AND2_X1 _25654_ (.A1(_08103_),
    .A2(_08132_),
    .ZN(_08134_));
 AOI221_X1 _25655_ (.A(_08133_),
    .B1(_08083_),
    .B2(_07651_),
    .C1(\cs_registers_i.mhpmcounter[2][21] ),
    .C2(_08134_),
    .ZN(_01766_));
 OR2_X1 _25656_ (.A1(\cs_registers_i.mhpmcounter[2][22] ),
    .A2(_08045_),
    .ZN(_08135_));
 AND2_X1 _25657_ (.A1(\cs_registers_i.mhpmcounter[2][21] ),
    .A2(_08132_),
    .ZN(_08136_));
 AOI21_X1 _25658_ (.A(_08135_),
    .B1(_08136_),
    .B2(_08108_),
    .ZN(_08137_));
 AND2_X1 _25659_ (.A1(_08108_),
    .A2(_08136_),
    .ZN(_08138_));
 AOI221_X1 _25660_ (.A(_08137_),
    .B1(_08083_),
    .B2(_07656_),
    .C1(\cs_registers_i.mhpmcounter[2][22] ),
    .C2(_08138_),
    .ZN(_01767_));
 OR2_X1 _25661_ (.A1(_04759_),
    .A2(_08045_),
    .ZN(_08139_));
 AND2_X1 _25662_ (.A1(\cs_registers_i.mhpmcounter[2][21] ),
    .A2(\cs_registers_i.mhpmcounter[2][22] ),
    .ZN(_08140_));
 AND2_X1 _25663_ (.A1(_08132_),
    .A2(_08140_),
    .ZN(_08141_));
 AOI21_X1 _25664_ (.A(_08139_),
    .B1(_08141_),
    .B2(_08105_),
    .ZN(_08142_));
 AND2_X1 _25665_ (.A1(_08103_),
    .A2(_08141_),
    .ZN(_08143_));
 AOI221_X1 _25666_ (.A(_08142_),
    .B1(_08083_),
    .B2(_07669_),
    .C1(_04759_),
    .C2(_08143_),
    .ZN(_01768_));
 NAND2_X1 _25667_ (.A1(_04901_),
    .A2(_08055_),
    .ZN(_08144_));
 AND3_X1 _25668_ (.A1(_04759_),
    .A2(_08108_),
    .A3(_08141_),
    .ZN(_08145_));
 BUF_X2 _25669_ (.A(_08048_),
    .Z(_08146_));
 NAND2_X1 _25670_ (.A1(_04759_),
    .A2(_08141_),
    .ZN(_08147_));
 NOR4_X1 _25671_ (.A1(_04901_),
    .A2(_08146_),
    .A3(_08107_),
    .A4(_08147_),
    .ZN(_08148_));
 INV_X4 _25672_ (.A(_07676_),
    .ZN(_08149_));
 AOI21_X1 _25673_ (.A(_08148_),
    .B1(_08112_),
    .B2(_08149_),
    .ZN(_08150_));
 OAI22_X1 _25674_ (.A1(_08144_),
    .A2(_08145_),
    .B1(_08150_),
    .B2(_08114_),
    .ZN(_01769_));
 NOR2_X1 _25675_ (.A1(_07689_),
    .A2(_08055_),
    .ZN(_08151_));
 INV_X1 _25676_ (.A(\cs_registers_i.mhpmcounter[2][25] ),
    .ZN(_08152_));
 NAND2_X1 _25677_ (.A1(_08152_),
    .A2(_08055_),
    .ZN(_08153_));
 AND3_X1 _25678_ (.A1(_04759_),
    .A2(_04901_),
    .A3(_08141_),
    .ZN(_08154_));
 AOI21_X1 _25679_ (.A(_08153_),
    .B1(_08154_),
    .B2(_08105_),
    .ZN(_08155_));
 AND3_X1 _25680_ (.A1(\cs_registers_i.mhpmcounter[2][25] ),
    .A2(_08105_),
    .A3(_08154_),
    .ZN(_08156_));
 NOR3_X1 _25681_ (.A1(_08151_),
    .A2(_08155_),
    .A3(_08156_),
    .ZN(_01770_));
 INV_X1 _25682_ (.A(\cs_registers_i.mhpmcounter[2][26] ),
    .ZN(_08157_));
 NAND2_X1 _25683_ (.A1(_08157_),
    .A2(_08054_),
    .ZN(_08158_));
 NAND4_X2 _25684_ (.A1(_04759_),
    .A2(_04901_),
    .A3(_08132_),
    .A4(_08140_),
    .ZN(_08159_));
 NOR2_X1 _25685_ (.A1(_08152_),
    .A2(_08159_),
    .ZN(_08160_));
 AOI21_X1 _25686_ (.A(_08158_),
    .B1(_08160_),
    .B2(_08108_),
    .ZN(_08161_));
 NOR3_X2 _25687_ (.A1(_08152_),
    .A2(_08157_),
    .A3(_08159_),
    .ZN(_08162_));
 BUF_X4 _25688_ (.A(_07696_),
    .Z(_08163_));
 AOI221_X1 _25689_ (.A(_08161_),
    .B1(_08162_),
    .B2(_08108_),
    .C1(_08047_),
    .C2(_08163_),
    .ZN(_01771_));
 NAND2_X1 _25690_ (.A1(\cs_registers_i.mhpmcounter[2][27] ),
    .A2(_08055_),
    .ZN(_08164_));
 AND2_X1 _25691_ (.A1(_08105_),
    .A2(_08162_),
    .ZN(_08165_));
 INV_X1 _25692_ (.A(\cs_registers_i.mhpmcounter[2][27] ),
    .ZN(_08166_));
 NAND3_X1 _25693_ (.A1(_08166_),
    .A2(_08101_),
    .A3(_08162_),
    .ZN(_08167_));
 MUX2_X1 _25694_ (.A(_07708_),
    .B(_08167_),
    .S(_08125_),
    .Z(_08168_));
 OAI22_X1 _25695_ (.A1(_08164_),
    .A2(_08165_),
    .B1(_08168_),
    .B2(_08114_),
    .ZN(_01772_));
 NAND2_X1 _25696_ (.A1(_05067_),
    .A2(_08055_),
    .ZN(_08169_));
 NOR4_X2 _25697_ (.A1(_08152_),
    .A2(_08157_),
    .A3(_08166_),
    .A4(_08159_),
    .ZN(_08170_));
 AND2_X1 _25698_ (.A1(_08108_),
    .A2(_08170_),
    .ZN(_08171_));
 INV_X1 _25699_ (.A(_08170_),
    .ZN(_08172_));
 NOR4_X1 _25700_ (.A1(_05067_),
    .A2(_08146_),
    .A3(_08107_),
    .A4(_08172_),
    .ZN(_08173_));
 AOI21_X1 _25701_ (.A(_08173_),
    .B1(_08112_),
    .B2(_07718_),
    .ZN(_08174_));
 OAI22_X1 _25702_ (.A1(_08169_),
    .A2(_08171_),
    .B1(_08174_),
    .B2(_08114_),
    .ZN(_01773_));
 OR2_X1 _25703_ (.A1(_05143_),
    .A2(_08045_),
    .ZN(_08175_));
 AND2_X1 _25704_ (.A1(_05067_),
    .A2(_08170_),
    .ZN(_08176_));
 AOI21_X1 _25705_ (.A(_08175_),
    .B1(_08176_),
    .B2(_08105_),
    .ZN(_08177_));
 AND2_X1 _25706_ (.A1(_08103_),
    .A2(_08176_),
    .ZN(_08178_));
 AOI221_X1 _25707_ (.A(_08177_),
    .B1(_08083_),
    .B2(_07727_),
    .C1(_05143_),
    .C2(_08178_),
    .ZN(_01774_));
 NAND2_X1 _25708_ (.A1(_04756_),
    .A2(_08039_),
    .ZN(_08179_));
 OAI21_X1 _25709_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .B1(_07492_),
    .B2(_08179_),
    .ZN(_08180_));
 MUX2_X1 _25710_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .B(_07493_),
    .S(_08041_),
    .Z(_08181_));
 NAND2_X1 _25711_ (.A1(_15532_),
    .A2(_08038_),
    .ZN(_08182_));
 MUX2_X1 _25712_ (.A(_08180_),
    .B(_08181_),
    .S(_08182_),
    .Z(_01775_));
 NOR2_X1 _25713_ (.A1(\cs_registers_i.mhpmcounter[2][30] ),
    .A2(_08047_),
    .ZN(_08183_));
 NAND4_X1 _25714_ (.A1(_04901_),
    .A2(\cs_registers_i.mhpmcounter[2][25] ),
    .A3(\cs_registers_i.mhpmcounter[2][26] ),
    .A4(\cs_registers_i.mhpmcounter[2][27] ),
    .ZN(_08184_));
 NOR2_X1 _25715_ (.A1(_08147_),
    .A2(_08184_),
    .ZN(_08185_));
 NAND4_X1 _25716_ (.A1(_05067_),
    .A2(_05143_),
    .A3(_08099_),
    .A4(_08185_),
    .ZN(_08186_));
 NAND3_X1 _25717_ (.A1(_08024_),
    .A2(_08029_),
    .A3(_08036_),
    .ZN(_08187_));
 OAI21_X1 _25718_ (.A(_08183_),
    .B1(_08186_),
    .B2(_08187_),
    .ZN(_08188_));
 NAND4_X1 _25719_ (.A1(_05067_),
    .A2(_05143_),
    .A3(\cs_registers_i.mhpmcounter[2][30] ),
    .A4(_08185_),
    .ZN(_08189_));
 NOR2_X1 _25720_ (.A1(_08107_),
    .A2(_08189_),
    .ZN(_08190_));
 AOI22_X1 _25721_ (.A1(_07983_),
    .A2(_08041_),
    .B1(_08190_),
    .B2(_08038_),
    .ZN(_08191_));
 AND2_X1 _25722_ (.A1(_08188_),
    .A2(_08191_),
    .ZN(_01776_));
 OR2_X1 _25723_ (.A1(\cs_registers_i.mhpmcounter[2][31] ),
    .A2(_08045_),
    .ZN(_08192_));
 AND4_X1 _25724_ (.A1(_05067_),
    .A2(_05143_),
    .A3(\cs_registers_i.mhpmcounter[2][30] ),
    .A4(_08170_),
    .ZN(_08193_));
 AOI21_X1 _25725_ (.A(_08192_),
    .B1(_08193_),
    .B2(_08105_),
    .ZN(_08194_));
 AND2_X1 _25726_ (.A1(_08103_),
    .A2(_08193_),
    .ZN(_08195_));
 AOI221_X1 _25727_ (.A(_08194_),
    .B1(_08083_),
    .B2(_07748_),
    .C1(\cs_registers_i.mhpmcounter[2][31] ),
    .C2(_08195_),
    .ZN(_01777_));
 AND2_X1 _25728_ (.A1(\cs_registers_i.mhpmcounter[2][31] ),
    .A2(_08193_),
    .ZN(_08196_));
 NAND2_X1 _25729_ (.A1(_08099_),
    .A2(_08196_),
    .ZN(_08197_));
 NAND2_X1 _25730_ (.A1(_08129_),
    .A2(_08197_),
    .ZN(_08198_));
 NOR2_X1 _25731_ (.A1(_04560_),
    .A2(_08043_),
    .ZN(_08199_));
 OAI33_X1 _25732_ (.A1(_04558_),
    .A2(_07487_),
    .A3(_08028_),
    .B1(net378),
    .B2(_08050_),
    .B3(_08199_),
    .ZN(_08200_));
 BUF_X4 _25733_ (.A(_08200_),
    .Z(_08201_));
 AOI21_X1 _25734_ (.A(_05352_),
    .B1(_08198_),
    .B2(_08201_),
    .ZN(_08202_));
 CLKBUF_X3 _25735_ (.A(_08125_),
    .Z(_08203_));
 OR2_X1 _25736_ (.A1(_08146_),
    .A2(_08197_),
    .ZN(_08204_));
 INV_X1 _25737_ (.A(_05352_),
    .ZN(_08205_));
 OAI22_X1 _25738_ (.A1(_07483_),
    .A2(_08203_),
    .B1(_08204_),
    .B2(_08205_),
    .ZN(_08206_));
 BUF_X4 _25739_ (.A(_08201_),
    .Z(_08207_));
 AOI21_X1 _25740_ (.A(_08202_),
    .B1(_08206_),
    .B2(_08207_),
    .ZN(_01778_));
 BUF_X8 _25741_ (.A(_08201_),
    .Z(_08208_));
 CLKBUF_X3 _25742_ (.A(_08125_),
    .Z(_08209_));
 NAND2_X1 _25743_ (.A1(_08101_),
    .A2(_08196_),
    .ZN(_08210_));
 OAI21_X1 _25744_ (.A(_08209_),
    .B1(_08210_),
    .B2(_08205_),
    .ZN(_08211_));
 AOI21_X1 _25745_ (.A(\cs_registers_i.mhpmcounter[2][33] ),
    .B1(_08208_),
    .B2(_08211_),
    .ZN(_08212_));
 NAND2_X1 _25746_ (.A1(_05352_),
    .A2(\cs_registers_i.mhpmcounter[2][33] ),
    .ZN(_08213_));
 NOR2_X1 _25747_ (.A1(_08210_),
    .A2(_08213_),
    .ZN(_08214_));
 CLKBUF_X3 _25748_ (.A(_08044_),
    .Z(_08215_));
 MUX2_X1 _25749_ (.A(_07635_),
    .B(_08214_),
    .S(_08215_),
    .Z(_08216_));
 AOI21_X1 _25750_ (.A(_08212_),
    .B1(_08216_),
    .B2(_08207_),
    .ZN(_01779_));
 OAI21_X1 _25751_ (.A(_08209_),
    .B1(_08197_),
    .B2(_08213_),
    .ZN(_08217_));
 AOI21_X1 _25752_ (.A(\cs_registers_i.mhpmcounter[2][34] ),
    .B1(_08208_),
    .B2(_08217_),
    .ZN(_08218_));
 NAND3_X1 _25753_ (.A1(_05352_),
    .A2(\cs_registers_i.mhpmcounter[2][33] ),
    .A3(\cs_registers_i.mhpmcounter[2][34] ),
    .ZN(_08219_));
 OAI22_X1 _25754_ (.A1(_07493_),
    .A2(_08203_),
    .B1(_08204_),
    .B2(_08219_),
    .ZN(_08220_));
 AOI21_X1 _25755_ (.A(_08218_),
    .B1(_08220_),
    .B2(_08207_),
    .ZN(_01780_));
 OR2_X1 _25756_ (.A1(_08210_),
    .A2(_08219_),
    .ZN(_08221_));
 NAND2_X1 _25757_ (.A1(_08129_),
    .A2(_08221_),
    .ZN(_08222_));
 AOI21_X1 _25758_ (.A(_05483_),
    .B1(_08208_),
    .B2(_08222_),
    .ZN(_08223_));
 INV_X1 _25759_ (.A(_07791_),
    .ZN(_08224_));
 OR2_X1 _25760_ (.A1(_08146_),
    .A2(_08221_),
    .ZN(_08225_));
 INV_X1 _25761_ (.A(_05483_),
    .ZN(_08226_));
 OAI22_X1 _25762_ (.A1(_08224_),
    .A2(_08203_),
    .B1(_08225_),
    .B2(_08226_),
    .ZN(_08227_));
 AOI21_X1 _25763_ (.A(_08223_),
    .B1(_08227_),
    .B2(_08207_),
    .ZN(_01781_));
 OR2_X1 _25764_ (.A1(_08197_),
    .A2(_08219_),
    .ZN(_08228_));
 OAI21_X1 _25765_ (.A(_08209_),
    .B1(_08228_),
    .B2(_08226_),
    .ZN(_08229_));
 AOI21_X1 _25766_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B1(_08208_),
    .B2(_08229_),
    .ZN(_08230_));
 INV_X2 _25767_ (.A(_07800_),
    .ZN(_08231_));
 NAND2_X1 _25768_ (.A1(_05483_),
    .A2(\cs_registers_i.mhpmcounter[2][36] ),
    .ZN(_08232_));
 OR2_X1 _25769_ (.A1(_08048_),
    .A2(_08228_),
    .ZN(_08233_));
 OAI22_X1 _25770_ (.A1(_08231_),
    .A2(_08203_),
    .B1(_08232_),
    .B2(_08233_),
    .ZN(_08234_));
 AOI21_X1 _25771_ (.A(_08230_),
    .B1(_08234_),
    .B2(_08207_),
    .ZN(_01782_));
 OAI21_X1 _25772_ (.A(_08209_),
    .B1(_08221_),
    .B2(_08232_),
    .ZN(_08235_));
 AOI21_X1 _25773_ (.A(\cs_registers_i.mhpmcounter[2][37] ),
    .B1(_08208_),
    .B2(_08235_),
    .ZN(_08236_));
 CLKBUF_X3 _25774_ (.A(_08125_),
    .Z(_08237_));
 NAND3_X2 _25775_ (.A1(_05483_),
    .A2(\cs_registers_i.mhpmcounter[2][36] ),
    .A3(\cs_registers_i.mhpmcounter[2][37] ),
    .ZN(_08238_));
 OAI22_X1 _25776_ (.A1(_07810_),
    .A2(_08237_),
    .B1(_08225_),
    .B2(_08238_),
    .ZN(_08239_));
 AOI21_X1 _25777_ (.A(_08236_),
    .B1(_08239_),
    .B2(_08207_),
    .ZN(_01783_));
 CLKBUF_X3 _25778_ (.A(_08125_),
    .Z(_08240_));
 OAI21_X1 _25779_ (.A(_08240_),
    .B1(_08228_),
    .B2(_08238_),
    .ZN(_08241_));
 AOI21_X1 _25780_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .B1(_08208_),
    .B2(_08241_),
    .ZN(_08242_));
 INV_X1 _25781_ (.A(_07821_),
    .ZN(_08243_));
 INV_X1 _25782_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .ZN(_08244_));
 OR2_X1 _25783_ (.A1(_08244_),
    .A2(_08238_),
    .ZN(_08245_));
 OAI22_X1 _25784_ (.A1(_08243_),
    .A2(_08237_),
    .B1(_08233_),
    .B2(_08245_),
    .ZN(_08246_));
 AOI21_X1 _25785_ (.A(_08242_),
    .B1(_08246_),
    .B2(_08207_),
    .ZN(_01784_));
 BUF_X8 _25786_ (.A(_08201_),
    .Z(_08247_));
 OAI21_X1 _25787_ (.A(_08240_),
    .B1(_08221_),
    .B2(_08245_),
    .ZN(_08248_));
 AOI21_X1 _25788_ (.A(\cs_registers_i.mhpmcounter[2][39] ),
    .B1(_08247_),
    .B2(_08248_),
    .ZN(_08249_));
 INV_X1 _25789_ (.A(_07828_),
    .ZN(_08250_));
 NOR2_X1 _25790_ (.A1(_08244_),
    .A2(_08238_),
    .ZN(_08251_));
 NAND2_X1 _25791_ (.A1(\cs_registers_i.mhpmcounter[2][39] ),
    .A2(_08251_),
    .ZN(_08252_));
 OAI22_X1 _25792_ (.A1(_08250_),
    .A2(_08237_),
    .B1(_08225_),
    .B2(_08252_),
    .ZN(_08253_));
 AOI21_X1 _25793_ (.A(_08249_),
    .B1(_08253_),
    .B2(_08207_),
    .ZN(_01785_));
 OR2_X1 _25794_ (.A1(\cs_registers_i.mhpmcounter[2][3] ),
    .A2(_08045_),
    .ZN(_08254_));
 AOI21_X1 _25795_ (.A(_08254_),
    .B1(_08069_),
    .B2(_08037_),
    .ZN(_08255_));
 AOI221_X2 _25796_ (.A(_08255_),
    .B1(_08080_),
    .B2(_08038_),
    .C1(_07791_),
    .C2(_08041_),
    .ZN(_01786_));
 OAI21_X1 _25797_ (.A(_08240_),
    .B1(_08228_),
    .B2(_08252_),
    .ZN(_08256_));
 AOI21_X1 _25798_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .B1(_08247_),
    .B2(_08256_),
    .ZN(_08257_));
 NAND3_X1 _25799_ (.A1(\cs_registers_i.mhpmcounter[2][39] ),
    .A2(\cs_registers_i.mhpmcounter[2][40] ),
    .A3(_08251_),
    .ZN(_08258_));
 OAI22_X1 _25800_ (.A1(_07844_),
    .A2(_08237_),
    .B1(_08233_),
    .B2(_08258_),
    .ZN(_08259_));
 AOI21_X1 _25801_ (.A(_08257_),
    .B1(_08259_),
    .B2(_08207_),
    .ZN(_01787_));
 OR2_X2 _25802_ (.A1(_08221_),
    .A2(_08258_),
    .ZN(_08260_));
 NAND2_X1 _25803_ (.A1(_08129_),
    .A2(_08260_),
    .ZN(_08261_));
 AOI21_X1 _25804_ (.A(_05708_),
    .B1(_08247_),
    .B2(_08261_),
    .ZN(_08262_));
 OR2_X1 _25805_ (.A1(_08146_),
    .A2(_08260_),
    .ZN(_08263_));
 INV_X1 _25806_ (.A(_05708_),
    .ZN(_08264_));
 OAI22_X1 _25807_ (.A1(_07854_),
    .A2(_08237_),
    .B1(_08263_),
    .B2(_08264_),
    .ZN(_08265_));
 AOI21_X1 _25808_ (.A(_08262_),
    .B1(_08265_),
    .B2(_08207_),
    .ZN(_01788_));
 OR2_X2 _25809_ (.A1(_08228_),
    .A2(_08258_),
    .ZN(_08266_));
 OAI21_X1 _25810_ (.A(_08240_),
    .B1(_08266_),
    .B2(_08264_),
    .ZN(_08267_));
 AOI21_X1 _25811_ (.A(\cs_registers_i.mhpmcounter[2][42] ),
    .B1(_08247_),
    .B2(_08267_),
    .ZN(_08268_));
 NAND2_X1 _25812_ (.A1(_05708_),
    .A2(\cs_registers_i.mhpmcounter[2][42] ),
    .ZN(_08269_));
 NOR2_X1 _25813_ (.A1(_08266_),
    .A2(_08269_),
    .ZN(_08270_));
 MUX2_X1 _25814_ (.A(_07525_),
    .B(_08270_),
    .S(_08215_),
    .Z(_08271_));
 BUF_X4 _25815_ (.A(_08201_),
    .Z(_08272_));
 AOI21_X1 _25816_ (.A(_08268_),
    .B1(_08271_),
    .B2(_08272_),
    .ZN(_01789_));
 OAI21_X1 _25817_ (.A(_08240_),
    .B1(_08260_),
    .B2(_08269_),
    .ZN(_08273_));
 AOI21_X1 _25818_ (.A(\cs_registers_i.mhpmcounter[2][43] ),
    .B1(_08247_),
    .B2(_08273_),
    .ZN(_08274_));
 INV_X2 _25819_ (.A(_07535_),
    .ZN(_08275_));
 NAND3_X1 _25820_ (.A1(\cs_registers_i.mhpmcounter[2][43] ),
    .A2(_05708_),
    .A3(\cs_registers_i.mhpmcounter[2][42] ),
    .ZN(_08276_));
 OAI22_X1 _25821_ (.A1(_08275_),
    .A2(_08237_),
    .B1(_08263_),
    .B2(_08276_),
    .ZN(_08277_));
 AOI21_X1 _25822_ (.A(_08274_),
    .B1(_08277_),
    .B2(_08272_),
    .ZN(_01790_));
 OAI21_X1 _25823_ (.A(_08240_),
    .B1(_08266_),
    .B2(_08276_),
    .ZN(_08278_));
 AOI21_X1 _25824_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .B1(_08247_),
    .B2(_08278_),
    .ZN(_08279_));
 INV_X1 _25825_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .ZN(_08280_));
 NOR3_X1 _25826_ (.A1(_08280_),
    .A2(_08266_),
    .A3(_08276_),
    .ZN(_08281_));
 MUX2_X1 _25827_ (.A(_07554_),
    .B(_08281_),
    .S(_08215_),
    .Z(_08282_));
 AOI21_X1 _25828_ (.A(_08279_),
    .B1(_08282_),
    .B2(_08272_),
    .ZN(_01791_));
 OR2_X1 _25829_ (.A1(_08280_),
    .A2(_08276_),
    .ZN(_08283_));
 OAI21_X1 _25830_ (.A(_08240_),
    .B1(_08260_),
    .B2(_08283_),
    .ZN(_08284_));
 AOI21_X1 _25831_ (.A(\cs_registers_i.mhpmcounter[2][45] ),
    .B1(_08247_),
    .B2(_08284_),
    .ZN(_08285_));
 INV_X1 _25832_ (.A(\cs_registers_i.mhpmcounter[2][45] ),
    .ZN(_08286_));
 OR2_X1 _25833_ (.A1(_08286_),
    .A2(_08283_),
    .ZN(_08287_));
 OAI22_X1 _25834_ (.A1(_07569_),
    .A2(_08237_),
    .B1(_08263_),
    .B2(_08287_),
    .ZN(_08288_));
 AOI21_X1 _25835_ (.A(_08285_),
    .B1(_08288_),
    .B2(_08272_),
    .ZN(_01792_));
 INV_X1 _25836_ (.A(_05914_),
    .ZN(_08289_));
 NOR2_X1 _25837_ (.A1(_08266_),
    .A2(_08287_),
    .ZN(_08290_));
 OAI21_X1 _25838_ (.A(_08208_),
    .B1(_08290_),
    .B2(_08112_),
    .ZN(_08291_));
 NAND3_X1 _25839_ (.A1(_05914_),
    .A2(_08215_),
    .A3(_08290_),
    .ZN(_08292_));
 OAI21_X1 _25840_ (.A(_08292_),
    .B1(_08237_),
    .B2(_07579_),
    .ZN(_08293_));
 AOI22_X1 _25841_ (.A1(_08289_),
    .A2(_08291_),
    .B1(_08293_),
    .B2(_08208_),
    .ZN(_01793_));
 NOR2_X1 _25842_ (.A1(_08260_),
    .A2(_08287_),
    .ZN(_08294_));
 NAND2_X1 _25843_ (.A1(_05914_),
    .A2(_08294_),
    .ZN(_08295_));
 NAND2_X1 _25844_ (.A1(_08129_),
    .A2(_08295_),
    .ZN(_08296_));
 AOI21_X1 _25845_ (.A(_05967_),
    .B1(_08247_),
    .B2(_08296_),
    .ZN(_08297_));
 NAND4_X1 _25846_ (.A1(_05914_),
    .A2(_05967_),
    .A3(_08209_),
    .A4(_08294_),
    .ZN(_08298_));
 INV_X2 _25847_ (.A(_07585_),
    .ZN(_08299_));
 OAI21_X1 _25848_ (.A(_08298_),
    .B1(_08203_),
    .B2(_08299_),
    .ZN(_08300_));
 AOI21_X1 _25849_ (.A(_08297_),
    .B1(_08300_),
    .B2(_08272_),
    .ZN(_01794_));
 NAND3_X1 _25850_ (.A1(_05914_),
    .A2(_05967_),
    .A3(_08290_),
    .ZN(_08301_));
 NAND2_X1 _25851_ (.A1(_08129_),
    .A2(_08301_),
    .ZN(_08302_));
 AOI21_X1 _25852_ (.A(\cs_registers_i.mhpmcounter[2][48] ),
    .B1(_08247_),
    .B2(_08302_),
    .ZN(_08303_));
 INV_X1 _25853_ (.A(\cs_registers_i.mhpmcounter[2][48] ),
    .ZN(_08304_));
 NOR2_X1 _25854_ (.A1(_08304_),
    .A2(_08301_),
    .ZN(_08305_));
 NAND2_X1 _25855_ (.A1(_08129_),
    .A2(_08305_),
    .ZN(_08306_));
 OAI21_X1 _25856_ (.A(_08306_),
    .B1(_08203_),
    .B2(_07600_),
    .ZN(_08307_));
 AOI21_X1 _25857_ (.A(_08303_),
    .B1(_08307_),
    .B2(_08272_),
    .ZN(_01795_));
 INV_X1 _25858_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .ZN(_08308_));
 NAND3_X1 _25859_ (.A1(_05914_),
    .A2(_05967_),
    .A3(\cs_registers_i.mhpmcounter[2][48] ),
    .ZN(_08309_));
 NOR3_X2 _25860_ (.A1(_08260_),
    .A2(_08287_),
    .A3(_08309_),
    .ZN(_08310_));
 OAI21_X1 _25861_ (.A(_08208_),
    .B1(_08310_),
    .B2(_08112_),
    .ZN(_08311_));
 BUF_X4 _25862_ (.A(_07605_),
    .Z(_08312_));
 NAND2_X1 _25863_ (.A1(_08312_),
    .A2(_08112_),
    .ZN(_08313_));
 NAND2_X2 _25864_ (.A1(\cs_registers_i.mhpmcounter[2][49] ),
    .A2(_08310_),
    .ZN(_08314_));
 OAI21_X1 _25865_ (.A(_08313_),
    .B1(_08314_),
    .B2(_08112_),
    .ZN(_08315_));
 AOI22_X1 _25866_ (.A1(_08308_),
    .A2(_08311_),
    .B1(_08315_),
    .B2(_08208_),
    .ZN(_01796_));
 NOR2_X1 _25867_ (.A1(_08231_),
    .A2(_08055_),
    .ZN(_08316_));
 OR2_X1 _25868_ (.A1(_05538_),
    .A2(_08046_),
    .ZN(_08317_));
 AOI21_X1 _25869_ (.A(_08317_),
    .B1(_08060_),
    .B2(_08038_),
    .ZN(_08318_));
 AND3_X1 _25870_ (.A1(_05538_),
    .A2(_08052_),
    .A3(_08060_),
    .ZN(_08319_));
 NOR3_X1 _25871_ (.A1(_08316_),
    .A2(_08318_),
    .A3(_08319_),
    .ZN(_01797_));
 NAND2_X2 _25872_ (.A1(\cs_registers_i.mhpmcounter[2][49] ),
    .A2(_08305_),
    .ZN(_08320_));
 NAND2_X1 _25873_ (.A1(_08129_),
    .A2(_08320_),
    .ZN(_08321_));
 AOI21_X1 _25874_ (.A(_06092_),
    .B1(_08247_),
    .B2(_08321_),
    .ZN(_08322_));
 NOR2_X1 _25875_ (.A1(_08146_),
    .A2(_08320_),
    .ZN(_08323_));
 AOI22_X1 _25876_ (.A1(_07616_),
    .A2(_08112_),
    .B1(_08323_),
    .B2(_06092_),
    .ZN(_08324_));
 INV_X1 _25877_ (.A(_08324_),
    .ZN(_08325_));
 AOI21_X1 _25878_ (.A(_08322_),
    .B1(_08325_),
    .B2(_08272_),
    .ZN(_01798_));
 BUF_X8 _25879_ (.A(_08201_),
    .Z(_08326_));
 INV_X1 _25880_ (.A(_06092_),
    .ZN(_08327_));
 OAI21_X1 _25881_ (.A(_08240_),
    .B1(_08314_),
    .B2(_08327_),
    .ZN(_08328_));
 AOI21_X1 _25882_ (.A(\cs_registers_i.mhpmcounter[2][51] ),
    .B1(_08326_),
    .B2(_08328_),
    .ZN(_08329_));
 NAND2_X1 _25883_ (.A1(_06092_),
    .A2(\cs_registers_i.mhpmcounter[2][51] ),
    .ZN(_08330_));
 NOR2_X1 _25884_ (.A1(_08314_),
    .A2(_08330_),
    .ZN(_08331_));
 MUX2_X1 _25885_ (.A(_07624_),
    .B(_08331_),
    .S(_08215_),
    .Z(_08332_));
 AOI21_X1 _25886_ (.A(_08329_),
    .B1(_08332_),
    .B2(_08272_),
    .ZN(_01799_));
 OAI21_X1 _25887_ (.A(_08240_),
    .B1(_08320_),
    .B2(_08330_),
    .ZN(_08333_));
 AOI21_X1 _25888_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .B1(_08326_),
    .B2(_08333_),
    .ZN(_08334_));
 NAND3_X1 _25889_ (.A1(_06092_),
    .A2(\cs_registers_i.mhpmcounter[2][51] ),
    .A3(\cs_registers_i.mhpmcounter[2][52] ),
    .ZN(_08335_));
 INV_X1 _25890_ (.A(_08335_),
    .ZN(_08336_));
 AOI22_X1 _25891_ (.A1(_07640_),
    .A2(_08112_),
    .B1(_08323_),
    .B2(_08336_),
    .ZN(_08337_));
 INV_X1 _25892_ (.A(_08337_),
    .ZN(_08338_));
 AOI21_X1 _25893_ (.A(_08334_),
    .B1(_08338_),
    .B2(_08272_),
    .ZN(_01800_));
 NOR2_X1 _25894_ (.A1(_08314_),
    .A2(_08335_),
    .ZN(_08339_));
 OR2_X1 _25895_ (.A1(_08146_),
    .A2(_08339_),
    .ZN(_08340_));
 AOI21_X1 _25896_ (.A(_06194_),
    .B1(_08326_),
    .B2(_08340_),
    .ZN(_08341_));
 NAND3_X1 _25897_ (.A1(_06194_),
    .A2(_08129_),
    .A3(_08339_),
    .ZN(_08342_));
 INV_X2 _25898_ (.A(_07651_),
    .ZN(_08343_));
 OAI21_X1 _25899_ (.A(_08342_),
    .B1(_08203_),
    .B2(_08343_),
    .ZN(_08344_));
 AOI21_X1 _25900_ (.A(_08341_),
    .B1(_08344_),
    .B2(_08272_),
    .ZN(_01801_));
 INV_X1 _25901_ (.A(_06194_),
    .ZN(_08345_));
 OAI33_X1 _25902_ (.A1(_07511_),
    .A2(_07487_),
    .A3(_08028_),
    .B1(_08320_),
    .B2(_08335_),
    .B3(_08345_),
    .ZN(_08346_));
 AOI21_X1 _25903_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .B1(_08326_),
    .B2(_08346_),
    .ZN(_08347_));
 NAND3_X1 _25904_ (.A1(_06194_),
    .A2(\cs_registers_i.mhpmcounter[2][54] ),
    .A3(_08336_),
    .ZN(_08348_));
 NOR2_X1 _25905_ (.A1(_08320_),
    .A2(_08348_),
    .ZN(_08349_));
 MUX2_X1 _25906_ (.A(_07657_),
    .B(_08349_),
    .S(_08215_),
    .Z(_08350_));
 BUF_X4 _25907_ (.A(_08201_),
    .Z(_08351_));
 AOI21_X1 _25908_ (.A(_08347_),
    .B1(_08350_),
    .B2(_08351_),
    .ZN(_01802_));
 OR2_X1 _25909_ (.A1(_08314_),
    .A2(_08348_),
    .ZN(_08352_));
 NAND2_X1 _25910_ (.A1(_08129_),
    .A2(_08352_),
    .ZN(_08353_));
 AOI21_X1 _25911_ (.A(_04754_),
    .B1(_08326_),
    .B2(_08353_),
    .ZN(_08354_));
 INV_X2 _25912_ (.A(_07669_),
    .ZN(_08355_));
 OR2_X1 _25913_ (.A1(_08146_),
    .A2(_08352_),
    .ZN(_08356_));
 INV_X1 _25914_ (.A(_04754_),
    .ZN(_08357_));
 OAI22_X1 _25915_ (.A1(_08355_),
    .A2(_08237_),
    .B1(_08356_),
    .B2(_08357_),
    .ZN(_08358_));
 AOI21_X1 _25916_ (.A(_08354_),
    .B1(_08358_),
    .B2(_08351_),
    .ZN(_01803_));
 NAND2_X1 _25917_ (.A1(_04754_),
    .A2(_08349_),
    .ZN(_08359_));
 NAND2_X1 _25918_ (.A1(_08209_),
    .A2(_08359_),
    .ZN(_08360_));
 AOI21_X1 _25919_ (.A(_04899_),
    .B1(_08326_),
    .B2(_08360_),
    .ZN(_08361_));
 NAND4_X1 _25920_ (.A1(_04754_),
    .A2(_04899_),
    .A3(_08209_),
    .A4(_08349_),
    .ZN(_08362_));
 OAI21_X1 _25921_ (.A(_08362_),
    .B1(_08203_),
    .B2(_08149_),
    .ZN(_08363_));
 AOI21_X1 _25922_ (.A(_08361_),
    .B1(_08363_),
    .B2(_08351_),
    .ZN(_01804_));
 NAND2_X1 _25923_ (.A1(_04754_),
    .A2(_04899_),
    .ZN(_08364_));
 OAI21_X1 _25924_ (.A(_08240_),
    .B1(_08352_),
    .B2(_08364_),
    .ZN(_08365_));
 AOI21_X1 _25925_ (.A(\cs_registers_i.mhpmcounter[2][57] ),
    .B1(_08326_),
    .B2(_08365_),
    .ZN(_08366_));
 NAND3_X1 _25926_ (.A1(_04754_),
    .A2(_04899_),
    .A3(\cs_registers_i.mhpmcounter[2][57] ),
    .ZN(_08367_));
 OAI22_X1 _25927_ (.A1(_07689_),
    .A2(_08237_),
    .B1(_08356_),
    .B2(_08367_),
    .ZN(_08368_));
 AOI21_X1 _25928_ (.A(_08366_),
    .B1(_08368_),
    .B2(_08351_),
    .ZN(_01805_));
 OR3_X2 _25929_ (.A1(_08320_),
    .A2(_08348_),
    .A3(_08367_),
    .ZN(_08369_));
 NAND2_X1 _25930_ (.A1(_08209_),
    .A2(_08369_),
    .ZN(_08370_));
 AOI21_X1 _25931_ (.A(_05029_),
    .B1(_08326_),
    .B2(_08370_),
    .ZN(_08371_));
 INV_X1 _25932_ (.A(_05029_),
    .ZN(_08372_));
 NOR3_X1 _25933_ (.A1(_08372_),
    .A2(_08146_),
    .A3(_08369_),
    .ZN(_08373_));
 AOI21_X1 _25934_ (.A(_08373_),
    .B1(_08112_),
    .B2(_08163_),
    .ZN(_08374_));
 INV_X1 _25935_ (.A(_08374_),
    .ZN(_08375_));
 AOI21_X1 _25936_ (.A(_08371_),
    .B1(_08375_),
    .B2(_08351_),
    .ZN(_01806_));
 OR2_X1 _25937_ (.A1(_08352_),
    .A2(_08367_),
    .ZN(_08376_));
 OAI21_X1 _25938_ (.A(_08215_),
    .B1(_08376_),
    .B2(_08372_),
    .ZN(_08377_));
 AOI21_X1 _25939_ (.A(_04781_),
    .B1(_08326_),
    .B2(_08377_),
    .ZN(_08378_));
 NAND2_X1 _25940_ (.A1(_05029_),
    .A2(_04781_),
    .ZN(_08379_));
 NOR2_X1 _25941_ (.A1(_08376_),
    .A2(_08379_),
    .ZN(_08380_));
 MUX2_X1 _25942_ (.A(_07708_),
    .B(_08380_),
    .S(_08125_),
    .Z(_08381_));
 AOI21_X1 _25943_ (.A(_08378_),
    .B1(_08381_),
    .B2(_08351_),
    .ZN(_01807_));
 NAND2_X1 _25944_ (.A1(_08061_),
    .A2(_08080_),
    .ZN(_08382_));
 OAI22_X1 _25945_ (.A1(_07810_),
    .A2(_08179_),
    .B1(_08382_),
    .B2(_08187_),
    .ZN(_08383_));
 NAND3_X1 _25946_ (.A1(_05538_),
    .A2(_08052_),
    .A3(_08080_),
    .ZN(_08384_));
 NOR2_X1 _25947_ (.A1(\cs_registers_i.mhpmcounter[2][5] ),
    .A2(_08047_),
    .ZN(_08385_));
 AOI21_X1 _25948_ (.A(_08383_),
    .B1(_08384_),
    .B2(_08385_),
    .ZN(_01808_));
 OAI21_X1 _25949_ (.A(_08215_),
    .B1(_08369_),
    .B2(_08379_),
    .ZN(_08386_));
 AOI21_X1 _25950_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .B1(_08326_),
    .B2(_08386_),
    .ZN(_08387_));
 NAND3_X1 _25951_ (.A1(_05029_),
    .A2(_04781_),
    .A3(\cs_registers_i.mhpmcounter[2][60] ),
    .ZN(_08388_));
 OR3_X1 _25952_ (.A1(_08146_),
    .A2(_08369_),
    .A3(_08388_),
    .ZN(_08389_));
 OAI21_X1 _25953_ (.A(_08389_),
    .B1(_08203_),
    .B2(_07718_),
    .ZN(_08390_));
 AOI21_X1 _25954_ (.A(_08387_),
    .B1(_08390_),
    .B2(_08351_),
    .ZN(_01809_));
 OAI21_X1 _25955_ (.A(_08215_),
    .B1(_08376_),
    .B2(_08388_),
    .ZN(_08391_));
 AOI21_X1 _25956_ (.A(\cs_registers_i.mhpmcounter[2][61] ),
    .B1(_08201_),
    .B2(_08391_),
    .ZN(_08392_));
 NAND4_X2 _25957_ (.A1(_05029_),
    .A2(_04781_),
    .A3(\cs_registers_i.mhpmcounter[2][60] ),
    .A4(\cs_registers_i.mhpmcounter[2][61] ),
    .ZN(_08393_));
 NOR2_X1 _25958_ (.A1(_08376_),
    .A2(_08393_),
    .ZN(_08394_));
 MUX2_X1 _25959_ (.A(_07728_),
    .B(_08394_),
    .S(_08125_),
    .Z(_08395_));
 AOI21_X1 _25960_ (.A(_08392_),
    .B1(_08395_),
    .B2(_08351_),
    .ZN(_01810_));
 OAI21_X1 _25961_ (.A(_08215_),
    .B1(_08369_),
    .B2(_08393_),
    .ZN(_08396_));
 AOI21_X1 _25962_ (.A(_05188_),
    .B1(_08201_),
    .B2(_08396_),
    .ZN(_08397_));
 INV_X1 _25963_ (.A(_05188_),
    .ZN(_08398_));
 NOR3_X1 _25964_ (.A1(_08398_),
    .A2(_08369_),
    .A3(_08393_),
    .ZN(_08399_));
 MUX2_X1 _25965_ (.A(_07745_),
    .B(_08399_),
    .S(_08125_),
    .Z(_08400_));
 AOI21_X1 _25966_ (.A(_08397_),
    .B1(_08400_),
    .B2(_08351_),
    .ZN(_01811_));
 NAND2_X1 _25967_ (.A1(_05188_),
    .A2(_08394_),
    .ZN(_08401_));
 NAND2_X1 _25968_ (.A1(_08209_),
    .A2(_08401_),
    .ZN(_08402_));
 AOI21_X1 _25969_ (.A(\cs_registers_i.mhpmcounter[2][63] ),
    .B1(_08201_),
    .B2(_08402_),
    .ZN(_08403_));
 NAND4_X1 _25970_ (.A1(_05188_),
    .A2(\cs_registers_i.mhpmcounter[2][63] ),
    .A3(_08209_),
    .A4(_08394_),
    .ZN(_08404_));
 INV_X2 _25971_ (.A(_07748_),
    .ZN(_08405_));
 OAI21_X1 _25972_ (.A(_08404_),
    .B1(_08203_),
    .B2(_08405_),
    .ZN(_08406_));
 AOI21_X1 _25973_ (.A(_08403_),
    .B1(_08406_),
    .B2(_08351_),
    .ZN(_01812_));
 OR2_X1 _25974_ (.A1(_05607_),
    .A2(_08045_),
    .ZN(_08407_));
 AOI21_X1 _25975_ (.A(_08407_),
    .B1(_08062_),
    .B2(_08037_),
    .ZN(_08408_));
 AND3_X1 _25976_ (.A1(_08051_),
    .A2(_08060_),
    .A3(_08061_),
    .ZN(_08409_));
 AOI221_X2 _25977_ (.A(_08408_),
    .B1(_08083_),
    .B2(_07821_),
    .C1(_05607_),
    .C2(_08409_),
    .ZN(_01813_));
 NOR2_X1 _25978_ (.A1(\cs_registers_i.mhpmcounter[2][7] ),
    .A2(_08046_),
    .ZN(_08410_));
 AND4_X1 _25979_ (.A1(_05607_),
    .A2(_08029_),
    .A3(_08061_),
    .A4(_08080_),
    .ZN(_08411_));
 NAND3_X1 _25980_ (.A1(_08024_),
    .A2(_08036_),
    .A3(_08411_),
    .ZN(_08412_));
 MUX2_X1 _25981_ (.A(\cs_registers_i.mhpmcounter[2][7] ),
    .B(_08410_),
    .S(_08412_),
    .Z(_08413_));
 AOI21_X1 _25982_ (.A(_08413_),
    .B1(_08047_),
    .B2(_07828_),
    .ZN(_01814_));
 NOR2_X1 _25983_ (.A1(_07844_),
    .A2(_08054_),
    .ZN(_08414_));
 AND3_X1 _25984_ (.A1(_05607_),
    .A2(\cs_registers_i.mhpmcounter[2][7] ),
    .A3(_08061_),
    .ZN(_08415_));
 AND4_X1 _25985_ (.A1(\cs_registers_i.mhpmcounter[2][8] ),
    .A2(_08051_),
    .A3(_08060_),
    .A4(_08415_),
    .ZN(_08416_));
 NAND3_X1 _25986_ (.A1(_08052_),
    .A2(_08060_),
    .A3(_08415_),
    .ZN(_08417_));
 NOR2_X1 _25987_ (.A1(\cs_registers_i.mhpmcounter[2][8] ),
    .A2(_08083_),
    .ZN(_08418_));
 AOI211_X2 _25988_ (.A(_08414_),
    .B(_08416_),
    .C1(_08417_),
    .C2(_08418_),
    .ZN(_01815_));
 NAND2_X1 _25989_ (.A1(_07854_),
    .A2(_08047_),
    .ZN(_08419_));
 INV_X1 _25990_ (.A(\cs_registers_i.mhpmcounter[2][9] ),
    .ZN(_08420_));
 AND2_X1 _25991_ (.A1(\cs_registers_i.mhpmcounter[2][8] ),
    .A2(_08415_),
    .ZN(_08421_));
 NAND4_X1 _25992_ (.A1(_08420_),
    .A2(_08052_),
    .A3(_08080_),
    .A4(_08421_),
    .ZN(_08422_));
 AND3_X1 _25993_ (.A1(_08052_),
    .A2(_08080_),
    .A3(_08421_),
    .ZN(_08423_));
 NAND2_X1 _25994_ (.A1(\cs_registers_i.mhpmcounter[2][9] ),
    .A2(_08055_),
    .ZN(_08424_));
 OAI211_X2 _25995_ (.A(_08419_),
    .B(_08422_),
    .C1(_08423_),
    .C2(_08424_),
    .ZN(_01816_));
 OAI21_X1 _25996_ (.A(_06989_),
    .B1(_06291_),
    .B2(_03850_),
    .ZN(_08425_));
 OR4_X2 _25997_ (.A1(_03436_),
    .A2(_03954_),
    .A3(_06293_),
    .A4(_03890_),
    .ZN(_08426_));
 NOR2_X2 _25998_ (.A1(_11420_),
    .A2(_03890_),
    .ZN(_08427_));
 NAND2_X4 _25999_ (.A1(_03880_),
    .A2(_08427_),
    .ZN(_08428_));
 AND2_X2 _26000_ (.A1(_03873_),
    .A2(_08428_),
    .ZN(_08429_));
 AND3_X1 _26001_ (.A1(_08425_),
    .A2(_08426_),
    .A3(_08429_),
    .ZN(_08430_));
 MUX2_X1 _26002_ (.A(_03462_),
    .B(\cs_registers_i.mstack_d[0] ),
    .S(_03924_),
    .Z(_08431_));
 NOR2_X1 _26003_ (.A1(_03927_),
    .A2(_08431_),
    .ZN(_08432_));
 NOR2_X1 _26004_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(_06803_),
    .ZN(_08433_));
 OAI21_X1 _26005_ (.A(_08430_),
    .B1(_08432_),
    .B2(_08433_),
    .ZN(_01817_));
 MUX2_X1 _26006_ (.A(_03463_),
    .B(\cs_registers_i.mstack_d[1] ),
    .S(_03924_),
    .Z(_08434_));
 NOR2_X1 _26007_ (.A1(_03927_),
    .A2(_08434_),
    .ZN(_08435_));
 NOR2_X1 _26008_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(_06803_),
    .ZN(_08436_));
 OAI21_X1 _26009_ (.A(_08430_),
    .B1(_08435_),
    .B2(_08436_),
    .ZN(_01818_));
 NAND2_X4 _26010_ (.A1(_08426_),
    .A2(_08428_),
    .ZN(_08437_));
 CLKBUF_X3 _26011_ (.A(_08437_),
    .Z(_08438_));
 NAND2_X1 _26012_ (.A1(_03462_),
    .A2(_08438_),
    .ZN(_08439_));
 AND2_X1 _26013_ (.A1(_05198_),
    .A2(_07489_),
    .ZN(_08440_));
 CLKBUF_X3 _26014_ (.A(_08440_),
    .Z(_08441_));
 NAND3_X1 _26015_ (.A1(_07482_),
    .A2(_07635_),
    .A3(_08441_),
    .ZN(_08442_));
 OAI21_X1 _26016_ (.A(_08442_),
    .B1(_08441_),
    .B2(\cs_registers_i.dcsr_q[0] ),
    .ZN(_08443_));
 OAI21_X1 _26017_ (.A(_08439_),
    .B1(_08443_),
    .B2(_08438_),
    .ZN(_01819_));
 MUX2_X1 _26018_ (.A(\cs_registers_i.dcsr_q[11] ),
    .B(_08275_),
    .S(_08441_),
    .Z(_01820_));
 INV_X1 _26019_ (.A(_07554_),
    .ZN(_08444_));
 MUX2_X1 _26020_ (.A(\cs_registers_i.dcsr_q[12] ),
    .B(_08444_),
    .S(_08441_),
    .Z(_01821_));
 MUX2_X1 _26021_ (.A(\cs_registers_i.dcsr_q[13] ),
    .B(_07569_),
    .S(_08441_),
    .Z(_01822_));
 MUX2_X1 _26022_ (.A(\cs_registers_i.dcsr_q[15] ),
    .B(_08299_),
    .S(_08441_),
    .Z(_01823_));
 NAND2_X1 _26023_ (.A1(_03463_),
    .A2(_08438_),
    .ZN(_08445_));
 OAI21_X1 _26024_ (.A(_08442_),
    .B1(_08441_),
    .B2(\cs_registers_i.dcsr_q[1] ),
    .ZN(_08446_));
 OAI21_X1 _26025_ (.A(_08445_),
    .B1(_08446_),
    .B2(_08438_),
    .ZN(_01824_));
 MUX2_X1 _26026_ (.A(_03879_),
    .B(_07493_),
    .S(_08441_),
    .Z(_01825_));
 AND2_X1 _26027_ (.A1(_08426_),
    .A2(_08428_),
    .ZN(_08447_));
 CLKBUF_X3 _26028_ (.A(_08447_),
    .Z(_08448_));
 INV_X1 _26029_ (.A(\cs_registers_i.dcsr_q[6] ),
    .ZN(_08449_));
 AOI22_X1 _26030_ (.A1(_03879_),
    .A2(_08427_),
    .B1(_08448_),
    .B2(_08449_),
    .ZN(_01826_));
 AOI22_X1 _26031_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_08426_),
    .B1(_08427_),
    .B2(net69),
    .ZN(_08450_));
 AOI21_X1 _26032_ (.A(_08450_),
    .B1(_08427_),
    .B2(_03879_),
    .ZN(_01827_));
 INV_X1 _26033_ (.A(\cs_registers_i.dcsr_q[8] ),
    .ZN(_08451_));
 OAI22_X1 _26034_ (.A1(_01162_),
    .A2(_08428_),
    .B1(_08438_),
    .B2(_08451_),
    .ZN(_01828_));
 NAND2_X2 _26035_ (.A1(_03873_),
    .A2(_08428_),
    .ZN(_08452_));
 BUF_X4 _26036_ (.A(_08452_),
    .Z(_08453_));
 BUF_X4 _26037_ (.A(_08453_),
    .Z(_08454_));
 MUX2_X1 _26038_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(\cs_registers_i.pc_if_i[10] ),
    .S(_08454_),
    .Z(_08455_));
 NAND2_X1 _26039_ (.A1(_08438_),
    .A2(_08455_),
    .ZN(_08456_));
 NAND2_X4 _26040_ (.A1(_04968_),
    .A2(_07489_),
    .ZN(_08457_));
 CLKBUF_X3 _26041_ (.A(_08457_),
    .Z(_08458_));
 NAND2_X2 _26042_ (.A1(_08448_),
    .A2(_08457_),
    .ZN(_08459_));
 CLKBUF_X3 _26043_ (.A(_08459_),
    .Z(_08460_));
 INV_X1 _26044_ (.A(\cs_registers_i.csr_depc_o[10] ),
    .ZN(_08461_));
 OAI221_X1 _26045_ (.A(_08456_),
    .B1(_08458_),
    .B2(_07525_),
    .C1(_08460_),
    .C2(_08461_),
    .ZN(_01829_));
 MUX2_X1 _26046_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_07178_),
    .S(_08454_),
    .Z(_08462_));
 NAND2_X1 _26047_ (.A1(_08438_),
    .A2(_08462_),
    .ZN(_08463_));
 INV_X1 _26048_ (.A(\cs_registers_i.csr_depc_o[11] ),
    .ZN(_08464_));
 OAI221_X1 _26049_ (.A(_08463_),
    .B1(_08458_),
    .B2(_07535_),
    .C1(_08464_),
    .C2(_08460_),
    .ZN(_01830_));
 MUX2_X1 _26050_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(_07199_),
    .S(_08454_),
    .Z(_08465_));
 NAND2_X1 _26051_ (.A1(_08438_),
    .A2(_08465_),
    .ZN(_08466_));
 INV_X1 _26052_ (.A(\cs_registers_i.csr_depc_o[12] ),
    .ZN(_08467_));
 OAI221_X1 _26053_ (.A(_08466_),
    .B1(_08458_),
    .B2(_07554_),
    .C1(_08467_),
    .C2(_08460_),
    .ZN(_01831_));
 NOR3_X4 _26054_ (.A1(_04260_),
    .A2(_04539_),
    .A3(_07487_),
    .ZN(_08468_));
 MUX2_X1 _26055_ (.A(_12076_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .S(_08453_),
    .Z(_08469_));
 CLKBUF_X3 _26056_ (.A(_08437_),
    .Z(_08470_));
 AOI22_X1 _26057_ (.A1(_07569_),
    .A2(_08468_),
    .B1(_08469_),
    .B2(_08470_),
    .ZN(_08471_));
 INV_X1 _26058_ (.A(\cs_registers_i.csr_depc_o[13] ),
    .ZN(_08472_));
 OAI21_X1 _26059_ (.A(_08471_),
    .B1(_08460_),
    .B2(_08472_),
    .ZN(_01832_));
 NOR2_X1 _26060_ (.A1(_07213_),
    .A2(_08429_),
    .ZN(_08473_));
 AOI21_X2 _26061_ (.A(_08473_),
    .B1(_08429_),
    .B2(_12179_),
    .ZN(_08474_));
 NAND2_X1 _26062_ (.A1(_08470_),
    .A2(_08474_),
    .ZN(_08475_));
 BUF_X4 _26063_ (.A(_08457_),
    .Z(_08476_));
 OAI221_X1 _26064_ (.A(_08475_),
    .B1(_08476_),
    .B2(_07579_),
    .C1(\cs_registers_i.csr_depc_o[14] ),
    .C2(_08459_),
    .ZN(_08477_));
 INV_X1 _26065_ (.A(_08477_),
    .ZN(_01833_));
 MUX2_X1 _26066_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_07222_),
    .S(_08454_),
    .Z(_08478_));
 NAND2_X1 _26067_ (.A1(_08438_),
    .A2(_08478_),
    .ZN(_08479_));
 INV_X1 _26068_ (.A(\cs_registers_i.csr_depc_o[15] ),
    .ZN(_08480_));
 OAI221_X1 _26069_ (.A(_08479_),
    .B1(_08458_),
    .B2(_07585_),
    .C1(_08480_),
    .C2(_08460_),
    .ZN(_01834_));
 NOR2_X1 _26070_ (.A1(_12352_),
    .A2(_08453_),
    .ZN(_08481_));
 AOI21_X2 _26071_ (.A(_08481_),
    .B1(_08454_),
    .B2(\cs_registers_i.pc_if_i[16] ),
    .ZN(_08482_));
 NOR2_X1 _26072_ (.A1(_08448_),
    .A2(_08482_),
    .ZN(_08483_));
 NOR2_X2 _26073_ (.A1(_08437_),
    .A2(_08468_),
    .ZN(_08484_));
 AOI221_X1 _26074_ (.A(_08483_),
    .B1(_08468_),
    .B2(_07600_),
    .C1(\cs_registers_i.csr_depc_o[16] ),
    .C2(_08484_),
    .ZN(_08485_));
 INV_X1 _26075_ (.A(_08485_),
    .ZN(_01835_));
 MUX2_X1 _26076_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(\cs_registers_i.pc_if_i[17] ),
    .S(_08453_),
    .Z(_08486_));
 NAND2_X1 _26077_ (.A1(_08438_),
    .A2(_08486_),
    .ZN(_08487_));
 OAI221_X1 _26078_ (.A(_08487_),
    .B1(_08458_),
    .B2(_08312_),
    .C1(_06051_),
    .C2(_08460_),
    .ZN(_01836_));
 CLKBUF_X3 _26079_ (.A(_08437_),
    .Z(_08488_));
 MUX2_X2 _26080_ (.A(\cs_registers_i.pc_id_i[18] ),
    .B(_07235_),
    .S(_08454_),
    .Z(_08489_));
 NAND2_X1 _26081_ (.A1(_08488_),
    .A2(_08489_),
    .ZN(_08490_));
 CLKBUF_X3 _26082_ (.A(_08459_),
    .Z(_08491_));
 OAI221_X1 _26083_ (.A(_08490_),
    .B1(_08458_),
    .B2(_07616_),
    .C1(_06954_),
    .C2(_08491_),
    .ZN(_01837_));
 BUF_X4 _26084_ (.A(_08452_),
    .Z(_08492_));
 MUX2_X1 _26085_ (.A(_12590_),
    .B(_07241_),
    .S(_08492_),
    .Z(_08493_));
 NOR2_X1 _26086_ (.A1(_08448_),
    .A2(_08493_),
    .ZN(_08494_));
 INV_X1 _26087_ (.A(\cs_registers_i.csr_depc_o[19] ),
    .ZN(_08495_));
 AOI221_X1 _26088_ (.A(_08494_),
    .B1(_08468_),
    .B2(_07623_),
    .C1(_08495_),
    .C2(_08484_),
    .ZN(_01838_));
 MUX2_X1 _26089_ (.A(_03981_),
    .B(_10675_),
    .S(_08429_),
    .Z(_08496_));
 NAND2_X1 _26090_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(_08457_),
    .ZN(_08497_));
 OAI21_X1 _26091_ (.A(_08497_),
    .B1(_08457_),
    .B2(_07635_),
    .ZN(_08498_));
 MUX2_X1 _26092_ (.A(_08496_),
    .B(_08498_),
    .S(_08448_),
    .Z(_01839_));
 MUX2_X1 _26093_ (.A(_12685_),
    .B(_07249_),
    .S(_08453_),
    .Z(_08499_));
 NOR2_X1 _26094_ (.A1(_08448_),
    .A2(_08499_),
    .ZN(_08500_));
 INV_X1 _26095_ (.A(\cs_registers_i.csr_depc_o[20] ),
    .ZN(_08501_));
 AOI221_X1 _26096_ (.A(_08500_),
    .B1(_08468_),
    .B2(_07639_),
    .C1(_08501_),
    .C2(_08484_),
    .ZN(_01840_));
 MUX2_X2 _26097_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(\cs_registers_i.pc_if_i[21] ),
    .S(_08454_),
    .Z(_08502_));
 NAND2_X1 _26098_ (.A1(_08488_),
    .A2(_08502_),
    .ZN(_08503_));
 OAI221_X1 _26099_ (.A(_08503_),
    .B1(_08458_),
    .B2(_07651_),
    .C1(_07000_),
    .C2(_08491_),
    .ZN(_01841_));
 MUX2_X2 _26100_ (.A(\cs_registers_i.pc_id_i[22] ),
    .B(_07259_),
    .S(_08492_),
    .Z(_08504_));
 NAND2_X1 _26101_ (.A1(_08488_),
    .A2(_08504_),
    .ZN(_08505_));
 OAI221_X1 _26102_ (.A(_08505_),
    .B1(_08458_),
    .B2(_07657_),
    .C1(_04540_),
    .C2(_08491_),
    .ZN(_01842_));
 MUX2_X1 _26103_ (.A(_12935_),
    .B(_07263_),
    .S(_08492_),
    .Z(_08506_));
 NAND2_X1 _26104_ (.A1(_08488_),
    .A2(_08506_),
    .ZN(_08507_));
 INV_X1 _26105_ (.A(\cs_registers_i.csr_depc_o[23] ),
    .ZN(_08508_));
 OAI221_X1 _26106_ (.A(_08507_),
    .B1(_08458_),
    .B2(_07669_),
    .C1(_08508_),
    .C2(_08491_),
    .ZN(_01843_));
 MUX2_X2 _26107_ (.A(_13024_),
    .B(\cs_registers_i.pc_if_i[24] ),
    .S(_08492_),
    .Z(_08509_));
 NAND2_X1 _26108_ (.A1(_08488_),
    .A2(_08509_),
    .ZN(_08510_));
 INV_X1 _26109_ (.A(\cs_registers_i.csr_depc_o[24] ),
    .ZN(_08511_));
 OAI221_X1 _26110_ (.A(_08510_),
    .B1(_08458_),
    .B2(_07676_),
    .C1(_08511_),
    .C2(_08491_),
    .ZN(_01844_));
 MUX2_X1 _26111_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(\cs_registers_i.pc_if_i[25] ),
    .S(_08453_),
    .Z(_08512_));
 AOI22_X1 _26112_ (.A1(_07689_),
    .A2(_08468_),
    .B1(_08512_),
    .B2(_08470_),
    .ZN(_08513_));
 INV_X1 _26113_ (.A(\cs_registers_i.csr_depc_o[25] ),
    .ZN(_08514_));
 OAI21_X1 _26114_ (.A(_08513_),
    .B1(_08460_),
    .B2(_08514_),
    .ZN(_01845_));
 MUX2_X1 _26115_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(_07281_),
    .S(_08492_),
    .Z(_08515_));
 NAND2_X1 _26116_ (.A1(_08488_),
    .A2(_08515_),
    .ZN(_08516_));
 OAI221_X1 _26117_ (.A(_08516_),
    .B1(_08476_),
    .B2(_08163_),
    .C1(_05025_),
    .C2(_08491_),
    .ZN(_01846_));
 MUX2_X2 _26118_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(_07285_),
    .S(_08492_),
    .Z(_08517_));
 NAND2_X1 _26119_ (.A1(_08488_),
    .A2(_08517_),
    .ZN(_08518_));
 INV_X1 _26120_ (.A(\cs_registers_i.csr_depc_o[27] ),
    .ZN(_08519_));
 OAI221_X1 _26121_ (.A(_08518_),
    .B1(_08476_),
    .B2(_07709_),
    .C1(_08519_),
    .C2(_08491_),
    .ZN(_01847_));
 AND2_X1 _26122_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_08429_),
    .ZN(_08520_));
 AOI21_X2 _26123_ (.A(_08520_),
    .B1(_08454_),
    .B2(\cs_registers_i.pc_if_i[28] ),
    .ZN(_08521_));
 NOR2_X1 _26124_ (.A1(_08448_),
    .A2(_08521_),
    .ZN(_08522_));
 AOI221_X1 _26125_ (.A(_08522_),
    .B1(_08468_),
    .B2(_07718_),
    .C1(\cs_registers_i.csr_depc_o[28] ),
    .C2(_08484_),
    .ZN(_08523_));
 INV_X1 _26126_ (.A(_08523_),
    .ZN(_01848_));
 MUX2_X2 _26127_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(\cs_registers_i.pc_if_i[29] ),
    .S(_08492_),
    .Z(_08524_));
 NAND2_X1 _26128_ (.A1(_08488_),
    .A2(_08524_),
    .ZN(_08525_));
 INV_X1 _26129_ (.A(\cs_registers_i.csr_depc_o[29] ),
    .ZN(_08526_));
 OAI221_X1 _26130_ (.A(_08525_),
    .B1(_08476_),
    .B2(_07728_),
    .C1(_08526_),
    .C2(_08491_),
    .ZN(_01849_));
 MUX2_X1 _26131_ (.A(_15352_),
    .B(_00012_),
    .S(_08429_),
    .Z(_08527_));
 OAI22_X1 _26132_ (.A1(_07492_),
    .A2(_08457_),
    .B1(_08527_),
    .B2(_08448_),
    .ZN(_08528_));
 AOI21_X1 _26133_ (.A(_08528_),
    .B1(_08484_),
    .B2(\cs_registers_i.csr_depc_o[2] ),
    .ZN(_08529_));
 INV_X1 _26134_ (.A(_08529_),
    .ZN(_01850_));
 MUX2_X1 _26135_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(\cs_registers_i.pc_if_i[30] ),
    .S(_08492_),
    .Z(_08530_));
 NAND2_X1 _26136_ (.A1(_08488_),
    .A2(_08530_),
    .ZN(_08531_));
 INV_X1 _26137_ (.A(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_08532_));
 OAI221_X1 _26138_ (.A(_08531_),
    .B1(_08476_),
    .B2(_07983_),
    .C1(_08532_),
    .C2(_08491_),
    .ZN(_01851_));
 MUX2_X1 _26139_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(\cs_registers_i.pc_if_i[31] ),
    .S(_08453_),
    .Z(_08533_));
 NAND2_X1 _26140_ (.A1(_08488_),
    .A2(_08533_),
    .ZN(_08534_));
 INV_X1 _26141_ (.A(\cs_registers_i.csr_depc_o[31] ),
    .ZN(_08535_));
 OAI221_X1 _26142_ (.A(_08534_),
    .B1(_08476_),
    .B2(_07748_),
    .C1(_08535_),
    .C2(_08491_),
    .ZN(_01852_));
 MUX2_X1 _26143_ (.A(_11517_),
    .B(_07181_),
    .S(_08453_),
    .Z(_08536_));
 NAND2_X1 _26144_ (.A1(_08470_),
    .A2(_08536_),
    .ZN(_08537_));
 INV_X1 _26145_ (.A(\cs_registers_i.csr_depc_o[3] ),
    .ZN(_08538_));
 OAI221_X1 _26146_ (.A(_08537_),
    .B1(_08476_),
    .B2(_07791_),
    .C1(_08538_),
    .C2(_08459_),
    .ZN(_01853_));
 MUX2_X1 _26147_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(_07186_),
    .S(_08454_),
    .Z(_08539_));
 NAND2_X1 _26148_ (.A1(_08470_),
    .A2(_08539_),
    .ZN(_08540_));
 INV_X1 _26149_ (.A(\cs_registers_i.csr_depc_o[4] ),
    .ZN(_08541_));
 OAI221_X1 _26150_ (.A(_08540_),
    .B1(_08476_),
    .B2(_07800_),
    .C1(_08541_),
    .C2(_08459_),
    .ZN(_01854_));
 MUX2_X1 _26151_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_07187_),
    .S(_08454_),
    .Z(_08542_));
 AOI22_X1 _26152_ (.A1(_07810_),
    .A2(_08468_),
    .B1(_08542_),
    .B2(_08470_),
    .ZN(_08543_));
 INV_X1 _26153_ (.A(\cs_registers_i.csr_depc_o[5] ),
    .ZN(_08544_));
 OAI21_X1 _26154_ (.A(_08543_),
    .B1(_08460_),
    .B2(_08544_),
    .ZN(_01855_));
 MUX2_X1 _26155_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(\cs_registers_i.pc_if_i[6] ),
    .S(_08492_),
    .Z(_08545_));
 NAND2_X1 _26156_ (.A1(_08470_),
    .A2(_08545_),
    .ZN(_08546_));
 INV_X1 _26157_ (.A(\cs_registers_i.csr_depc_o[6] ),
    .ZN(_08547_));
 OAI221_X1 _26158_ (.A(_08546_),
    .B1(_08476_),
    .B2(_07821_),
    .C1(_08547_),
    .C2(_08459_),
    .ZN(_01856_));
 MUX2_X1 _26159_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_07185_),
    .S(_08492_),
    .Z(_08548_));
 NAND2_X1 _26160_ (.A1(_08470_),
    .A2(_08548_),
    .ZN(_08549_));
 INV_X1 _26161_ (.A(\cs_registers_i.csr_depc_o[7] ),
    .ZN(_08550_));
 OAI221_X1 _26162_ (.A(_08549_),
    .B1(_08476_),
    .B2(_07828_),
    .C1(_08550_),
    .C2(_08459_),
    .ZN(_01857_));
 MUX2_X1 _26163_ (.A(_11788_),
    .B(\cs_registers_i.pc_if_i[8] ),
    .S(_08453_),
    .Z(_08551_));
 AOI22_X1 _26164_ (.A1(_07844_),
    .A2(_08468_),
    .B1(_08551_),
    .B2(_08470_),
    .ZN(_08552_));
 INV_X1 _26165_ (.A(\cs_registers_i.csr_depc_o[8] ),
    .ZN(_08553_));
 OAI21_X1 _26166_ (.A(_08552_),
    .B1(_08460_),
    .B2(_08553_),
    .ZN(_01858_));
 MUX2_X1 _26167_ (.A(_11826_),
    .B(_07184_),
    .S(_08453_),
    .Z(_08554_));
 AOI22_X1 _26168_ (.A1(_07854_),
    .A2(_08468_),
    .B1(_08554_),
    .B2(_08470_),
    .ZN(_08555_));
 INV_X1 _26169_ (.A(\cs_registers_i.csr_depc_o[9] ),
    .ZN(_08556_));
 OAI21_X1 _26170_ (.A(_08555_),
    .B1(_08460_),
    .B2(_08556_),
    .ZN(_01859_));
 NAND2_X2 _26171_ (.A1(_04511_),
    .A2(_07489_),
    .ZN(_08557_));
 BUF_X4 _26172_ (.A(_08557_),
    .Z(_08558_));
 MUX2_X1 _26173_ (.A(_07483_),
    .B(\cs_registers_i.dscratch0_q[0] ),
    .S(_08558_),
    .Z(_01860_));
 CLKBUF_X3 _26174_ (.A(_08557_),
    .Z(_08559_));
 NAND2_X1 _26175_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(_08559_),
    .ZN(_08560_));
 CLKBUF_X3 _26176_ (.A(_08557_),
    .Z(_08561_));
 OAI21_X1 _26177_ (.A(_08560_),
    .B1(_08561_),
    .B2(_07525_),
    .ZN(_01861_));
 MUX2_X1 _26178_ (.A(_08275_),
    .B(\cs_registers_i.dscratch0_q[11] ),
    .S(_08558_),
    .Z(_01862_));
 MUX2_X1 _26179_ (.A(_08444_),
    .B(\cs_registers_i.dscratch0_q[12] ),
    .S(_08558_),
    .Z(_01863_));
 MUX2_X1 _26180_ (.A(_07569_),
    .B(\cs_registers_i.dscratch0_q[13] ),
    .S(_08558_),
    .Z(_01864_));
 MUX2_X1 _26181_ (.A(_07579_),
    .B(\cs_registers_i.dscratch0_q[14] ),
    .S(_08558_),
    .Z(_01865_));
 MUX2_X1 _26182_ (.A(_08299_),
    .B(\cs_registers_i.dscratch0_q[15] ),
    .S(_08558_),
    .Z(_01866_));
 MUX2_X1 _26183_ (.A(_07600_),
    .B(\cs_registers_i.dscratch0_q[16] ),
    .S(_08558_),
    .Z(_01867_));
 NAND2_X1 _26184_ (.A1(\cs_registers_i.dscratch0_q[17] ),
    .A2(_08559_),
    .ZN(_08562_));
 OAI21_X1 _26185_ (.A(_08562_),
    .B1(_08561_),
    .B2(_08312_),
    .ZN(_01868_));
 MUX2_X1 _26186_ (.A(_07914_),
    .B(\cs_registers_i.dscratch0_q[18] ),
    .S(_08558_),
    .Z(_01869_));
 NAND2_X1 _26187_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(_08559_),
    .ZN(_08563_));
 OAI21_X1 _26188_ (.A(_08563_),
    .B1(_08561_),
    .B2(_07624_),
    .ZN(_01870_));
 NAND2_X1 _26189_ (.A1(\cs_registers_i.dscratch0_q[1] ),
    .A2(_08559_),
    .ZN(_08564_));
 OAI21_X1 _26190_ (.A(_08564_),
    .B1(_08561_),
    .B2(_07635_),
    .ZN(_01871_));
 NAND2_X1 _26191_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_08559_),
    .ZN(_08565_));
 OAI21_X1 _26192_ (.A(_08565_),
    .B1(_08561_),
    .B2(_07640_),
    .ZN(_01872_));
 MUX2_X1 _26193_ (.A(_08343_),
    .B(\cs_registers_i.dscratch0_q[21] ),
    .S(_08558_),
    .Z(_01873_));
 NAND2_X1 _26194_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_08559_),
    .ZN(_08566_));
 OAI21_X1 _26195_ (.A(_08566_),
    .B1(_08561_),
    .B2(_07657_),
    .ZN(_01874_));
 MUX2_X1 _26196_ (.A(_08355_),
    .B(\cs_registers_i.dscratch0_q[23] ),
    .S(_08558_),
    .Z(_01875_));
 BUF_X4 _26197_ (.A(_08557_),
    .Z(_08567_));
 MUX2_X1 _26198_ (.A(_08149_),
    .B(\cs_registers_i.dscratch0_q[24] ),
    .S(_08567_),
    .Z(_01876_));
 MUX2_X1 _26199_ (.A(_07689_),
    .B(\cs_registers_i.dscratch0_q[25] ),
    .S(_08567_),
    .Z(_01877_));
 NAND2_X1 _26200_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(_08559_),
    .ZN(_08568_));
 OAI21_X1 _26201_ (.A(_08568_),
    .B1(_08561_),
    .B2(_08163_),
    .ZN(_01878_));
 NAND2_X1 _26202_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_08559_),
    .ZN(_08569_));
 OAI21_X1 _26203_ (.A(_08569_),
    .B1(_08561_),
    .B2(_07709_),
    .ZN(_01879_));
 MUX2_X1 _26204_ (.A(_07718_),
    .B(\cs_registers_i.dscratch0_q[28] ),
    .S(_08567_),
    .Z(_01880_));
 NAND2_X1 _26205_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(_08559_),
    .ZN(_08570_));
 OAI21_X1 _26206_ (.A(_08570_),
    .B1(_08561_),
    .B2(_07728_),
    .ZN(_01881_));
 MUX2_X1 _26207_ (.A(_07493_),
    .B(\cs_registers_i.dscratch0_q[2] ),
    .S(_08567_),
    .Z(_01882_));
 NAND2_X1 _26208_ (.A1(\cs_registers_i.dscratch0_q[30] ),
    .A2(_08559_),
    .ZN(_08571_));
 OAI21_X1 _26209_ (.A(_08571_),
    .B1(_08561_),
    .B2(_07983_),
    .ZN(_01883_));
 MUX2_X1 _26210_ (.A(_08405_),
    .B(\cs_registers_i.dscratch0_q[31] ),
    .S(_08567_),
    .Z(_01884_));
 MUX2_X1 _26211_ (.A(_08224_),
    .B(\cs_registers_i.dscratch0_q[3] ),
    .S(_08567_),
    .Z(_01885_));
 MUX2_X1 _26212_ (.A(_08231_),
    .B(\cs_registers_i.dscratch0_q[4] ),
    .S(_08567_),
    .Z(_01886_));
 MUX2_X1 _26213_ (.A(_07810_),
    .B(\cs_registers_i.dscratch0_q[5] ),
    .S(_08567_),
    .Z(_01887_));
 MUX2_X1 _26214_ (.A(_08243_),
    .B(\cs_registers_i.dscratch0_q[6] ),
    .S(_08567_),
    .Z(_01888_));
 MUX2_X1 _26215_ (.A(_08250_),
    .B(\cs_registers_i.dscratch0_q[7] ),
    .S(_08567_),
    .Z(_01889_));
 MUX2_X1 _26216_ (.A(_07844_),
    .B(\cs_registers_i.dscratch0_q[8] ),
    .S(_08557_),
    .Z(_01890_));
 MUX2_X1 _26217_ (.A(_07854_),
    .B(\cs_registers_i.dscratch0_q[9] ),
    .S(_08557_),
    .Z(_01891_));
 NAND2_X2 _26218_ (.A1(_04530_),
    .A2(_07489_),
    .ZN(_08572_));
 BUF_X4 _26219_ (.A(_08572_),
    .Z(_08573_));
 MUX2_X1 _26220_ (.A(_07483_),
    .B(\cs_registers_i.dscratch1_q[0] ),
    .S(_08573_),
    .Z(_01892_));
 CLKBUF_X3 _26221_ (.A(_08572_),
    .Z(_08574_));
 NAND2_X1 _26222_ (.A1(\cs_registers_i.dscratch1_q[10] ),
    .A2(_08574_),
    .ZN(_08575_));
 CLKBUF_X3 _26223_ (.A(_08572_),
    .Z(_08576_));
 OAI21_X1 _26224_ (.A(_08575_),
    .B1(_08576_),
    .B2(_07525_),
    .ZN(_01893_));
 MUX2_X1 _26225_ (.A(_08275_),
    .B(\cs_registers_i.dscratch1_q[11] ),
    .S(_08573_),
    .Z(_01894_));
 MUX2_X1 _26226_ (.A(_08444_),
    .B(\cs_registers_i.dscratch1_q[12] ),
    .S(_08573_),
    .Z(_01895_));
 MUX2_X1 _26227_ (.A(_07569_),
    .B(\cs_registers_i.dscratch1_q[13] ),
    .S(_08573_),
    .Z(_01896_));
 MUX2_X1 _26228_ (.A(_07579_),
    .B(\cs_registers_i.dscratch1_q[14] ),
    .S(_08573_),
    .Z(_01897_));
 MUX2_X1 _26229_ (.A(_08299_),
    .B(\cs_registers_i.dscratch1_q[15] ),
    .S(_08573_),
    .Z(_01898_));
 MUX2_X1 _26230_ (.A(_07600_),
    .B(\cs_registers_i.dscratch1_q[16] ),
    .S(_08573_),
    .Z(_01899_));
 NAND2_X1 _26231_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_08574_),
    .ZN(_08577_));
 OAI21_X1 _26232_ (.A(_08577_),
    .B1(_08576_),
    .B2(_08312_),
    .ZN(_01900_));
 MUX2_X1 _26233_ (.A(_07914_),
    .B(\cs_registers_i.dscratch1_q[18] ),
    .S(_08573_),
    .Z(_01901_));
 NAND2_X1 _26234_ (.A1(\cs_registers_i.dscratch1_q[19] ),
    .A2(_08574_),
    .ZN(_08578_));
 OAI21_X1 _26235_ (.A(_08578_),
    .B1(_08576_),
    .B2(_07624_),
    .ZN(_01902_));
 NAND2_X1 _26236_ (.A1(\cs_registers_i.dscratch1_q[1] ),
    .A2(_08574_),
    .ZN(_08579_));
 OAI21_X1 _26237_ (.A(_08579_),
    .B1(_08576_),
    .B2(_07635_),
    .ZN(_01903_));
 NAND2_X1 _26238_ (.A1(\cs_registers_i.dscratch1_q[20] ),
    .A2(_08574_),
    .ZN(_08580_));
 OAI21_X1 _26239_ (.A(_08580_),
    .B1(_08576_),
    .B2(_07640_),
    .ZN(_01904_));
 MUX2_X1 _26240_ (.A(_08343_),
    .B(\cs_registers_i.dscratch1_q[21] ),
    .S(_08573_),
    .Z(_01905_));
 NAND2_X1 _26241_ (.A1(\cs_registers_i.dscratch1_q[22] ),
    .A2(_08574_),
    .ZN(_08581_));
 OAI21_X1 _26242_ (.A(_08581_),
    .B1(_08576_),
    .B2(_07657_),
    .ZN(_01906_));
 MUX2_X1 _26243_ (.A(_08355_),
    .B(\cs_registers_i.dscratch1_q[23] ),
    .S(_08573_),
    .Z(_01907_));
 BUF_X4 _26244_ (.A(_08572_),
    .Z(_08582_));
 MUX2_X1 _26245_ (.A(_08149_),
    .B(\cs_registers_i.dscratch1_q[24] ),
    .S(_08582_),
    .Z(_01908_));
 MUX2_X1 _26246_ (.A(_07689_),
    .B(\cs_registers_i.dscratch1_q[25] ),
    .S(_08582_),
    .Z(_01909_));
 NAND2_X1 _26247_ (.A1(\cs_registers_i.dscratch1_q[26] ),
    .A2(_08574_),
    .ZN(_08583_));
 OAI21_X1 _26248_ (.A(_08583_),
    .B1(_08576_),
    .B2(_08163_),
    .ZN(_01910_));
 NAND2_X1 _26249_ (.A1(\cs_registers_i.dscratch1_q[27] ),
    .A2(_08574_),
    .ZN(_08584_));
 OAI21_X1 _26250_ (.A(_08584_),
    .B1(_08576_),
    .B2(_07709_),
    .ZN(_01911_));
 MUX2_X1 _26251_ (.A(_07718_),
    .B(\cs_registers_i.dscratch1_q[28] ),
    .S(_08582_),
    .Z(_01912_));
 NAND2_X1 _26252_ (.A1(\cs_registers_i.dscratch1_q[29] ),
    .A2(_08574_),
    .ZN(_08585_));
 OAI21_X1 _26253_ (.A(_08585_),
    .B1(_08576_),
    .B2(_07728_),
    .ZN(_01913_));
 MUX2_X1 _26254_ (.A(_07493_),
    .B(\cs_registers_i.dscratch1_q[2] ),
    .S(_08582_),
    .Z(_01914_));
 NAND2_X1 _26255_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_08574_),
    .ZN(_08586_));
 OAI21_X1 _26256_ (.A(_08586_),
    .B1(_08576_),
    .B2(_07983_),
    .ZN(_01915_));
 MUX2_X1 _26257_ (.A(_08405_),
    .B(\cs_registers_i.dscratch1_q[31] ),
    .S(_08582_),
    .Z(_01916_));
 MUX2_X1 _26258_ (.A(_08224_),
    .B(\cs_registers_i.dscratch1_q[3] ),
    .S(_08582_),
    .Z(_01917_));
 MUX2_X1 _26259_ (.A(_08231_),
    .B(\cs_registers_i.dscratch1_q[4] ),
    .S(_08582_),
    .Z(_01918_));
 MUX2_X1 _26260_ (.A(_07810_),
    .B(\cs_registers_i.dscratch1_q[5] ),
    .S(_08582_),
    .Z(_01919_));
 MUX2_X1 _26261_ (.A(_08243_),
    .B(\cs_registers_i.dscratch1_q[6] ),
    .S(_08582_),
    .Z(_01920_));
 MUX2_X1 _26262_ (.A(_08250_),
    .B(\cs_registers_i.dscratch1_q[7] ),
    .S(_08582_),
    .Z(_01921_));
 MUX2_X1 _26263_ (.A(_07844_),
    .B(\cs_registers_i.dscratch1_q[8] ),
    .S(_08572_),
    .Z(_01922_));
 MUX2_X1 _26264_ (.A(_07854_),
    .B(\cs_registers_i.dscratch1_q[9] ),
    .S(_08572_),
    .Z(_01923_));
 NOR3_X4 _26265_ (.A1(_03918_),
    .A2(_03894_),
    .A3(_03921_),
    .ZN(_08587_));
 BUF_X4 _26266_ (.A(_08587_),
    .Z(_08588_));
 NAND2_X1 _26267_ (.A1(\cs_registers_i.mstack_cause_q[0] ),
    .A2(_08588_),
    .ZN(_08589_));
 NAND2_X4 _26268_ (.A1(_03870_),
    .A2(_06797_),
    .ZN(_08590_));
 NOR2_X2 _26269_ (.A1(_08430_),
    .A2(_08437_),
    .ZN(_08591_));
 NAND2_X4 _26270_ (.A1(_03478_),
    .A2(_08591_),
    .ZN(_08592_));
 NAND2_X1 _26271_ (.A1(_08590_),
    .A2(_08592_),
    .ZN(_08593_));
 BUF_X4 _26272_ (.A(_08593_),
    .Z(_08594_));
 BUF_X4 _26273_ (.A(_08592_),
    .Z(_08595_));
 CLKBUF_X3 _26274_ (.A(_08595_),
    .Z(_08596_));
 CLKBUF_X3 _26275_ (.A(_06989_),
    .Z(_08597_));
 BUF_X4 _26276_ (.A(_03843_),
    .Z(_08598_));
 BUF_X4 _26277_ (.A(_08598_),
    .Z(_08599_));
 INV_X1 _26278_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .ZN(_08600_));
 BUF_X4 _26279_ (.A(_03842_),
    .Z(_08601_));
 NAND4_X4 _26280_ (.A1(_08600_),
    .A2(_08601_),
    .A3(_03610_),
    .A4(_03837_),
    .ZN(_08602_));
 BUF_X4 _26281_ (.A(_08602_),
    .Z(_08603_));
 INV_X1 _26282_ (.A(_08601_),
    .ZN(_08604_));
 NOR2_X1 _26283_ (.A1(_11935_),
    .A2(_08604_),
    .ZN(_08605_));
 NAND4_X1 _26284_ (.A1(_03435_),
    .A2(_03464_),
    .A3(_03609_),
    .A4(_08605_),
    .ZN(_08606_));
 OAI21_X1 _26285_ (.A(_08606_),
    .B1(_06291_),
    .B2(_03849_),
    .ZN(_08607_));
 NAND2_X1 _26286_ (.A1(_08601_),
    .A2(_08607_),
    .ZN(_08608_));
 NAND3_X1 _26287_ (.A1(_08599_),
    .A2(_08603_),
    .A3(_08608_),
    .ZN(_08609_));
 AOI21_X1 _26288_ (.A(_03920_),
    .B1(_08597_),
    .B2(_08609_),
    .ZN(_08610_));
 OAI221_X1 _26289_ (.A(_08589_),
    .B1(_08594_),
    .B2(_07482_),
    .C1(_08596_),
    .C2(_08610_),
    .ZN(_08611_));
 NAND2_X2 _26290_ (.A1(_03844_),
    .A2(_08591_),
    .ZN(_08612_));
 NAND2_X2 _26291_ (.A1(_08612_),
    .A2(_08590_),
    .ZN(_08613_));
 AOI21_X4 _26292_ (.A(_08613_),
    .B1(_07489_),
    .B2(_05228_),
    .ZN(_08614_));
 MUX2_X1 _26293_ (.A(_08611_),
    .B(\cs_registers_i.mcause_q[0] ),
    .S(_08614_),
    .Z(_01924_));
 OR2_X2 _26294_ (.A1(_08430_),
    .A2(_08437_),
    .ZN(_08615_));
 NOR2_X4 _26295_ (.A1(_03477_),
    .A2(_08615_),
    .ZN(_08616_));
 NOR2_X4 _26296_ (.A1(_08587_),
    .A2(_08616_),
    .ZN(_08617_));
 BUF_X4 _26297_ (.A(_08617_),
    .Z(_08618_));
 AND2_X1 _26298_ (.A1(_07634_),
    .A2(_08618_),
    .ZN(_08619_));
 BUF_X4 _26299_ (.A(_08616_),
    .Z(_08620_));
 NAND2_X2 _26300_ (.A1(_03461_),
    .A2(_03891_),
    .ZN(_08621_));
 NOR2_X1 _26301_ (.A1(_03607_),
    .A2(_08621_),
    .ZN(_08622_));
 NAND3_X1 _26302_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(_08600_),
    .A3(_08598_),
    .ZN(_08623_));
 NOR2_X1 _26303_ (.A1(_03609_),
    .A2(_08623_),
    .ZN(_08624_));
 NOR2_X1 _26304_ (.A1(_03849_),
    .A2(_03852_),
    .ZN(_08625_));
 AOI21_X1 _26305_ (.A(_08624_),
    .B1(_08625_),
    .B2(_03609_),
    .ZN(_08626_));
 NAND3_X1 _26306_ (.A1(_08601_),
    .A2(_08606_),
    .A3(_08626_),
    .ZN(_08627_));
 NAND2_X1 _26307_ (.A1(_08622_),
    .A2(_08627_),
    .ZN(_08628_));
 NAND3_X1 _26308_ (.A1(_03949_),
    .A2(_08620_),
    .A3(_08628_),
    .ZN(_08629_));
 OAI21_X1 _26309_ (.A(_08629_),
    .B1(_08590_),
    .B2(\cs_registers_i.mstack_cause_q[1] ),
    .ZN(_08630_));
 NOR2_X1 _26310_ (.A1(_08619_),
    .A2(_08630_),
    .ZN(_08631_));
 MUX2_X1 _26311_ (.A(_08631_),
    .B(\cs_registers_i.mcause_q[1] ),
    .S(_08614_),
    .Z(_01925_));
 NAND2_X1 _26312_ (.A1(\cs_registers_i.mcause_q[2] ),
    .A2(_08614_),
    .ZN(_08632_));
 BUF_X4 _26313_ (.A(_08620_),
    .Z(_08633_));
 NAND2_X1 _26314_ (.A1(_08598_),
    .A2(_06989_),
    .ZN(_08634_));
 OAI221_X1 _26315_ (.A(_08633_),
    .B1(_08603_),
    .B2(_08634_),
    .C1(_06802_),
    .C2(_03873_),
    .ZN(_08635_));
 BUF_X4 _26316_ (.A(_08593_),
    .Z(_08636_));
 INV_X1 _26317_ (.A(_08587_),
    .ZN(_08637_));
 OAI221_X1 _26318_ (.A(_08635_),
    .B1(_08636_),
    .B2(_07493_),
    .C1(\cs_registers_i.mstack_cause_q[2] ),
    .C2(_08637_),
    .ZN(_08638_));
 OAI21_X1 _26319_ (.A(_08632_),
    .B1(_08638_),
    .B2(_08614_),
    .ZN(_01926_));
 AND3_X1 _26320_ (.A1(_03609_),
    .A2(_08605_),
    .A3(_08622_),
    .ZN(_08639_));
 NOR3_X1 _26321_ (.A1(_06811_),
    .A2(_08592_),
    .A3(_08639_),
    .ZN(_08640_));
 INV_X1 _26322_ (.A(\cs_registers_i.mstack_cause_q[3] ),
    .ZN(_08641_));
 AOI221_X1 _26323_ (.A(_08640_),
    .B1(_08617_),
    .B2(_07791_),
    .C1(_08641_),
    .C2(_08587_),
    .ZN(_08642_));
 MUX2_X1 _26324_ (.A(_08642_),
    .B(\cs_registers_i.mcause_q[3] ),
    .S(_08614_),
    .Z(_01927_));
 NAND2_X1 _26325_ (.A1(\cs_registers_i.mcause_q[4] ),
    .A2(_08614_),
    .ZN(_08643_));
 NAND2_X1 _26326_ (.A1(_07800_),
    .A2(_08618_),
    .ZN(_08644_));
 OAI221_X1 _26327_ (.A(_08644_),
    .B1(_08596_),
    .B2(_06844_),
    .C1(\cs_registers_i.mstack_cause_q[4] ),
    .C2(_08637_),
    .ZN(_08645_));
 OAI21_X1 _26328_ (.A(_08643_),
    .B1(_08645_),
    .B2(_08614_),
    .ZN(_01928_));
 INV_X1 _26329_ (.A(\cs_registers_i.mcause_q[5] ),
    .ZN(_08646_));
 CLKBUF_X3 _26330_ (.A(_08616_),
    .Z(_08647_));
 NOR3_X1 _26331_ (.A1(_07748_),
    .A2(_08588_),
    .A3(_08647_),
    .ZN(_08648_));
 AOI21_X1 _26332_ (.A(_08648_),
    .B1(_08588_),
    .B2(\cs_registers_i.mstack_cause_q[5] ),
    .ZN(_08649_));
 NOR2_X1 _26333_ (.A1(_03941_),
    .A2(_08614_),
    .ZN(_08650_));
 AOI22_X1 _26334_ (.A1(_08646_),
    .A2(_08614_),
    .B1(_08649_),
    .B2(_08650_),
    .ZN(_01929_));
 AOI21_X4 _26335_ (.A(_08613_),
    .B1(_07489_),
    .B2(_04544_),
    .ZN(_08651_));
 AOI22_X1 _26336_ (.A1(\cs_registers_i.mstack_epc_q[0] ),
    .A2(_08588_),
    .B1(_08651_),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_08652_));
 INV_X1 _26337_ (.A(_08652_),
    .ZN(_01930_));
 BUF_X4 _26338_ (.A(_08587_),
    .Z(_08653_));
 AOI22_X1 _26339_ (.A1(\cs_registers_i.mstack_epc_q[10] ),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08455_),
    .ZN(_08654_));
 OAI21_X1 _26340_ (.A(_08654_),
    .B1(_08636_),
    .B2(_07525_),
    .ZN(_08655_));
 NAND2_X1 _26341_ (.A1(_04544_),
    .A2(_07488_),
    .ZN(_08656_));
 NAND3_X4 _26342_ (.A1(_08612_),
    .A2(_08590_),
    .A3(_08656_),
    .ZN(_08657_));
 BUF_X4 _26343_ (.A(_08657_),
    .Z(_08658_));
 MUX2_X1 _26344_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(_08655_),
    .S(_08658_),
    .Z(_01931_));
 AOI22_X1 _26345_ (.A1(\cs_registers_i.mstack_epc_q[11] ),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08462_),
    .ZN(_08659_));
 OAI21_X1 _26346_ (.A(_08659_),
    .B1(_08636_),
    .B2(_07535_),
    .ZN(_08660_));
 MUX2_X1 _26347_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(_08660_),
    .S(_08658_),
    .Z(_01932_));
 AOI22_X1 _26348_ (.A1(\cs_registers_i.mstack_epc_q[12] ),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08465_),
    .ZN(_08661_));
 OAI21_X1 _26349_ (.A(_08661_),
    .B1(_08636_),
    .B2(_07554_),
    .ZN(_08662_));
 MUX2_X1 _26350_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(_08662_),
    .S(_08658_),
    .Z(_01933_));
 CLKBUF_X3 _26351_ (.A(_08657_),
    .Z(_08663_));
 NOR2_X1 _26352_ (.A1(\cs_registers_i.csr_mepc_o[13] ),
    .A2(_08663_),
    .ZN(_08664_));
 AND2_X1 _26353_ (.A1(_08469_),
    .A2(_08616_),
    .ZN(_08665_));
 AOI221_X1 _26354_ (.A(_08665_),
    .B1(_08618_),
    .B2(_07568_),
    .C1(\cs_registers_i.mstack_epc_q[13] ),
    .C2(_08588_),
    .ZN(_08666_));
 AOI21_X1 _26355_ (.A(_08664_),
    .B1(_08666_),
    .B2(_08663_),
    .ZN(_01934_));
 NOR2_X1 _26356_ (.A1(\cs_registers_i.csr_mepc_o[14] ),
    .A2(_08663_),
    .ZN(_08667_));
 NOR2_X1 _26357_ (.A1(_08474_),
    .A2(_08592_),
    .ZN(_08668_));
 AOI221_X2 _26358_ (.A(_08668_),
    .B1(_08618_),
    .B2(_07579_),
    .C1(\cs_registers_i.mstack_epc_q[14] ),
    .C2(_08588_),
    .ZN(_08669_));
 AOI21_X1 _26359_ (.A(_08667_),
    .B1(_08669_),
    .B2(_08663_),
    .ZN(_01935_));
 AOI22_X1 _26360_ (.A1(\cs_registers_i.mstack_epc_q[15] ),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08478_),
    .ZN(_08670_));
 OAI21_X1 _26361_ (.A(_08670_),
    .B1(_08636_),
    .B2(_07585_),
    .ZN(_08671_));
 MUX2_X1 _26362_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(_08671_),
    .S(_08658_),
    .Z(_01936_));
 NOR2_X1 _26363_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_08663_),
    .ZN(_08672_));
 NOR2_X1 _26364_ (.A1(_08482_),
    .A2(_08592_),
    .ZN(_08673_));
 AOI221_X2 _26365_ (.A(_08673_),
    .B1(_08618_),
    .B2(_07600_),
    .C1(\cs_registers_i.mstack_epc_q[16] ),
    .C2(_08653_),
    .ZN(_08674_));
 AOI21_X1 _26366_ (.A(_08672_),
    .B1(_08674_),
    .B2(_08663_),
    .ZN(_01937_));
 AOI22_X1 _26367_ (.A1(\cs_registers_i.mstack_epc_q[17] ),
    .A2(_08587_),
    .B1(_08620_),
    .B2(_08486_),
    .ZN(_08675_));
 OAI21_X1 _26368_ (.A(_08675_),
    .B1(_08594_),
    .B2(_08312_),
    .ZN(_08676_));
 MUX2_X1 _26369_ (.A(_08676_),
    .B(\cs_registers_i.csr_mepc_o[17] ),
    .S(_08651_),
    .Z(_01938_));
 AOI22_X1 _26370_ (.A1(\cs_registers_i.mstack_epc_q[18] ),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08489_),
    .ZN(_08677_));
 OAI21_X1 _26371_ (.A(_08677_),
    .B1(_08636_),
    .B2(_07616_),
    .ZN(_08678_));
 MUX2_X1 _26372_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(_08678_),
    .S(_08658_),
    .Z(_01939_));
 CLKBUF_X3 _26373_ (.A(_08587_),
    .Z(_08679_));
 AOI22_X1 _26374_ (.A1(\cs_registers_i.mstack_epc_q[19] ),
    .A2(_08679_),
    .B1(_08647_),
    .B2(_08493_),
    .ZN(_08680_));
 OAI21_X1 _26375_ (.A(_08680_),
    .B1(_08636_),
    .B2(_07624_),
    .ZN(_08681_));
 MUX2_X1 _26376_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(_08681_),
    .S(_08658_),
    .Z(_01940_));
 OAI22_X1 _26377_ (.A1(\cs_registers_i.mstack_epc_q[1] ),
    .A2(_08590_),
    .B1(_08595_),
    .B2(_08496_),
    .ZN(_08682_));
 NOR2_X1 _26378_ (.A1(_08619_),
    .A2(_08682_),
    .ZN(_08683_));
 BUF_X4 _26379_ (.A(_08657_),
    .Z(_08684_));
 MUX2_X1 _26380_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(_08683_),
    .S(_08684_),
    .Z(_01941_));
 CLKBUF_X3 _26381_ (.A(_08616_),
    .Z(_08685_));
 AOI22_X1 _26382_ (.A1(\cs_registers_i.mstack_epc_q[20] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08499_),
    .ZN(_08686_));
 OAI21_X1 _26383_ (.A(_08686_),
    .B1(_08636_),
    .B2(_07640_),
    .ZN(_08687_));
 MUX2_X1 _26384_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(_08687_),
    .S(_08684_),
    .Z(_01942_));
 AOI22_X1 _26385_ (.A1(\cs_registers_i.mstack_epc_q[21] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08502_),
    .ZN(_08688_));
 OAI21_X1 _26386_ (.A(_08688_),
    .B1(_08636_),
    .B2(_07651_),
    .ZN(_08689_));
 MUX2_X1 _26387_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(_08689_),
    .S(_08684_),
    .Z(_01943_));
 AOI22_X1 _26388_ (.A1(\cs_registers_i.mstack_epc_q[22] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08504_),
    .ZN(_08690_));
 OAI21_X1 _26389_ (.A(_08690_),
    .B1(_08636_),
    .B2(_07657_),
    .ZN(_08691_));
 MUX2_X1 _26390_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(_08691_),
    .S(_08684_),
    .Z(_01944_));
 AOI22_X1 _26391_ (.A1(\cs_registers_i.mstack_epc_q[23] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08506_),
    .ZN(_08692_));
 OAI21_X1 _26392_ (.A(_08692_),
    .B1(_08594_),
    .B2(_07669_),
    .ZN(_08693_));
 MUX2_X1 _26393_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(_08693_),
    .S(_08684_),
    .Z(_01945_));
 AOI22_X1 _26394_ (.A1(\cs_registers_i.mstack_epc_q[24] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08509_),
    .ZN(_08694_));
 OAI21_X1 _26395_ (.A(_08694_),
    .B1(_08594_),
    .B2(_07676_),
    .ZN(_08695_));
 MUX2_X1 _26396_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(_08695_),
    .S(_08684_),
    .Z(_01946_));
 NOR2_X1 _26397_ (.A1(\cs_registers_i.csr_mepc_o[25] ),
    .A2(_08658_),
    .ZN(_08696_));
 AND2_X1 _26398_ (.A1(_08512_),
    .A2(_08616_),
    .ZN(_08697_));
 AOI221_X1 _26399_ (.A(_08697_),
    .B1(_08618_),
    .B2(_07688_),
    .C1(\cs_registers_i.mstack_epc_q[25] ),
    .C2(_08653_),
    .ZN(_08698_));
 AOI21_X1 _26400_ (.A(_08696_),
    .B1(_08698_),
    .B2(_08663_),
    .ZN(_01947_));
 AOI22_X1 _26401_ (.A1(\cs_registers_i.mstack_epc_q[26] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08515_),
    .ZN(_08699_));
 OAI21_X1 _26402_ (.A(_08699_),
    .B1(_08594_),
    .B2(_08163_),
    .ZN(_08700_));
 MUX2_X1 _26403_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(_08700_),
    .S(_08684_),
    .Z(_01948_));
 AOI22_X1 _26404_ (.A1(\cs_registers_i.mstack_epc_q[27] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08517_),
    .ZN(_08701_));
 OAI21_X1 _26405_ (.A(_08701_),
    .B1(_08594_),
    .B2(_07709_),
    .ZN(_08702_));
 MUX2_X1 _26406_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(_08702_),
    .S(_08684_),
    .Z(_01949_));
 NOR2_X1 _26407_ (.A1(\cs_registers_i.csr_mepc_o[28] ),
    .A2(_08658_),
    .ZN(_08703_));
 NOR2_X1 _26408_ (.A1(_08521_),
    .A2(_08592_),
    .ZN(_08704_));
 AOI221_X1 _26409_ (.A(_08704_),
    .B1(_08618_),
    .B2(_07717_),
    .C1(\cs_registers_i.mstack_epc_q[28] ),
    .C2(_08653_),
    .ZN(_08705_));
 AOI21_X1 _26410_ (.A(_08703_),
    .B1(_08705_),
    .B2(_08663_),
    .ZN(_01950_));
 AOI22_X1 _26411_ (.A1(\cs_registers_i.mstack_epc_q[29] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08524_),
    .ZN(_08706_));
 OAI21_X1 _26412_ (.A(_08706_),
    .B1(_08594_),
    .B2(_07728_),
    .ZN(_08707_));
 MUX2_X1 _26413_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(_08707_),
    .S(_08684_),
    .Z(_01951_));
 NOR2_X1 _26414_ (.A1(\cs_registers_i.mstack_epc_q[2] ),
    .A2(_08637_),
    .ZN(_08708_));
 AOI221_X1 _26415_ (.A(_08708_),
    .B1(_08620_),
    .B2(_08527_),
    .C1(_07492_),
    .C2(_08617_),
    .ZN(_08709_));
 MUX2_X1 _26416_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .B(_08709_),
    .S(_08684_),
    .Z(_01952_));
 AOI22_X1 _26417_ (.A1(\cs_registers_i.mstack_epc_q[30] ),
    .A2(_08679_),
    .B1(_08685_),
    .B2(_08530_),
    .ZN(_08710_));
 OAI21_X1 _26418_ (.A(_08710_),
    .B1(_08594_),
    .B2(_07983_),
    .ZN(_08711_));
 MUX2_X1 _26419_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(_08711_),
    .S(_08657_),
    .Z(_01953_));
 OAI22_X1 _26420_ (.A1(\cs_registers_i.mstack_epc_q[31] ),
    .A2(_08590_),
    .B1(_08595_),
    .B2(_08533_),
    .ZN(_08712_));
 AOI21_X1 _26421_ (.A(_08712_),
    .B1(_08618_),
    .B2(_07748_),
    .ZN(_08713_));
 MUX2_X1 _26422_ (.A(_08713_),
    .B(\cs_registers_i.csr_mepc_o[31] ),
    .S(_08651_),
    .Z(_01954_));
 OAI22_X1 _26423_ (.A1(\cs_registers_i.mstack_epc_q[3] ),
    .A2(_08590_),
    .B1(_08595_),
    .B2(_08536_),
    .ZN(_08714_));
 AOI21_X1 _26424_ (.A(_08714_),
    .B1(_08618_),
    .B2(_07791_),
    .ZN(_08715_));
 MUX2_X1 _26425_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(_08715_),
    .S(_08657_),
    .Z(_01955_));
 NAND2_X1 _26426_ (.A1(\cs_registers_i.csr_mepc_o[4] ),
    .A2(_08651_),
    .ZN(_08716_));
 OAI221_X1 _26427_ (.A(_08644_),
    .B1(_08596_),
    .B2(_08539_),
    .C1(\cs_registers_i.mstack_epc_q[4] ),
    .C2(_08637_),
    .ZN(_08717_));
 OAI21_X1 _26428_ (.A(_08716_),
    .B1(_08717_),
    .B2(_08651_),
    .ZN(_01956_));
 AOI22_X1 _26429_ (.A1(\cs_registers_i.mstack_epc_q[5] ),
    .A2(_08588_),
    .B1(_08647_),
    .B2(_08542_),
    .ZN(_08718_));
 NAND2_X1 _26430_ (.A1(_07810_),
    .A2(_08618_),
    .ZN(_08719_));
 AND3_X1 _26431_ (.A1(_08657_),
    .A2(_08718_),
    .A3(_08719_),
    .ZN(_08720_));
 AOI21_X1 _26432_ (.A(_08720_),
    .B1(_08651_),
    .B2(_06812_),
    .ZN(_01957_));
 AOI22_X1 _26433_ (.A1(\cs_registers_i.mstack_epc_q[6] ),
    .A2(_08587_),
    .B1(_08685_),
    .B2(_08545_),
    .ZN(_08721_));
 OAI21_X1 _26434_ (.A(_08721_),
    .B1(_08594_),
    .B2(_07821_),
    .ZN(_08722_));
 MUX2_X1 _26435_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(_08722_),
    .S(_08657_),
    .Z(_01958_));
 AOI22_X1 _26436_ (.A1(\cs_registers_i.mstack_epc_q[7] ),
    .A2(_08587_),
    .B1(_08620_),
    .B2(_08548_),
    .ZN(_08723_));
 OAI21_X1 _26437_ (.A(_08723_),
    .B1(_08594_),
    .B2(_07828_),
    .ZN(_08724_));
 MUX2_X1 _26438_ (.A(\cs_registers_i.csr_mepc_o[7] ),
    .B(_08724_),
    .S(_08657_),
    .Z(_01959_));
 NOR2_X1 _26439_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(_08658_),
    .ZN(_08725_));
 AND2_X1 _26440_ (.A1(_08551_),
    .A2(_08616_),
    .ZN(_08726_));
 AOI221_X1 _26441_ (.A(_08726_),
    .B1(_08617_),
    .B2(_07844_),
    .C1(\cs_registers_i.mstack_epc_q[8] ),
    .C2(_08653_),
    .ZN(_08727_));
 AOI21_X1 _26442_ (.A(_08725_),
    .B1(_08727_),
    .B2(_08663_),
    .ZN(_01960_));
 NOR2_X1 _26443_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_08658_),
    .ZN(_08728_));
 AND2_X1 _26444_ (.A1(_08554_),
    .A2(_08616_),
    .ZN(_08729_));
 AOI221_X2 _26445_ (.A(_08729_),
    .B1(_08617_),
    .B2(_07853_),
    .C1(\cs_registers_i.mstack_epc_q[9] ),
    .C2(_08653_),
    .ZN(_08730_));
 AOI21_X1 _26446_ (.A(_08728_),
    .B1(_08730_),
    .B2(_08663_),
    .ZN(_01961_));
 NAND2_X4 _26447_ (.A1(_04515_),
    .A2(_07489_),
    .ZN(_08731_));
 CLKBUF_X3 _26448_ (.A(_08731_),
    .Z(_08732_));
 MUX2_X1 _26449_ (.A(_07600_),
    .B(\cs_registers_i.mie_q[0] ),
    .S(_08732_),
    .Z(_01962_));
 CLKBUF_X3 _26450_ (.A(_08731_),
    .Z(_08733_));
 NAND2_X1 _26451_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(_08733_),
    .ZN(_08734_));
 OAI21_X1 _26452_ (.A(_08734_),
    .B1(_08733_),
    .B2(_08163_),
    .ZN(_01963_));
 NAND2_X1 _26453_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(_08733_),
    .ZN(_08735_));
 OAI21_X1 _26454_ (.A(_08735_),
    .B1(_08733_),
    .B2(_07709_),
    .ZN(_01964_));
 MUX2_X1 _26455_ (.A(_07718_),
    .B(\cs_registers_i.mie_q[12] ),
    .S(_08732_),
    .Z(_01965_));
 NAND2_X1 _26456_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(_08732_),
    .ZN(_08736_));
 OAI21_X1 _26457_ (.A(_08736_),
    .B1(_08733_),
    .B2(_07728_),
    .ZN(_01966_));
 NAND2_X1 _26458_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(_08732_),
    .ZN(_08737_));
 OAI21_X1 _26459_ (.A(_08737_),
    .B1(_08733_),
    .B2(_07983_),
    .ZN(_01967_));
 MUX2_X1 _26460_ (.A(_08275_),
    .B(\cs_registers_i.mie_q[15] ),
    .S(_08732_),
    .Z(_01968_));
 MUX2_X1 _26461_ (.A(_08250_),
    .B(\cs_registers_i.mie_q[16] ),
    .S(_08732_),
    .Z(_01969_));
 MUX2_X1 _26462_ (.A(_08224_),
    .B(\cs_registers_i.mie_q[17] ),
    .S(_08731_),
    .Z(_01970_));
 NAND2_X1 _26463_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(_08732_),
    .ZN(_08738_));
 OAI21_X1 _26464_ (.A(_08738_),
    .B1(_08733_),
    .B2(_08312_),
    .ZN(_01971_));
 MUX2_X1 _26465_ (.A(_07914_),
    .B(\cs_registers_i.mie_q[2] ),
    .S(_08731_),
    .Z(_01972_));
 NAND2_X1 _26466_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(_08732_),
    .ZN(_08739_));
 OAI21_X1 _26467_ (.A(_08739_),
    .B1(_08733_),
    .B2(_07624_),
    .ZN(_01973_));
 NAND2_X1 _26468_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(_08732_),
    .ZN(_08740_));
 OAI21_X1 _26469_ (.A(_08740_),
    .B1(_08733_),
    .B2(_07640_),
    .ZN(_01974_));
 MUX2_X1 _26470_ (.A(_08343_),
    .B(\cs_registers_i.mie_q[5] ),
    .S(_08731_),
    .Z(_01975_));
 NAND2_X1 _26471_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(_08732_),
    .ZN(_08741_));
 OAI21_X1 _26472_ (.A(_08741_),
    .B1(_08733_),
    .B2(_07657_),
    .ZN(_01976_));
 MUX2_X1 _26473_ (.A(_08355_),
    .B(\cs_registers_i.mie_q[7] ),
    .S(_08731_),
    .Z(_01977_));
 MUX2_X1 _26474_ (.A(_08149_),
    .B(\cs_registers_i.mie_q[8] ),
    .S(_08731_),
    .Z(_01978_));
 MUX2_X1 _26475_ (.A(_07689_),
    .B(\cs_registers_i.mie_q[9] ),
    .S(_08731_),
    .Z(_01979_));
 NAND2_X2 _26476_ (.A1(_04524_),
    .A2(_07489_),
    .ZN(_08742_));
 BUF_X4 _26477_ (.A(_08742_),
    .Z(_08743_));
 MUX2_X1 _26478_ (.A(_07483_),
    .B(\cs_registers_i.mscratch_q[0] ),
    .S(_08743_),
    .Z(_01980_));
 CLKBUF_X3 _26479_ (.A(_08742_),
    .Z(_08744_));
 NAND2_X1 _26480_ (.A1(\cs_registers_i.mscratch_q[10] ),
    .A2(_08744_),
    .ZN(_08745_));
 CLKBUF_X3 _26481_ (.A(_08742_),
    .Z(_08746_));
 OAI21_X1 _26482_ (.A(_08745_),
    .B1(_08746_),
    .B2(_07525_),
    .ZN(_01981_));
 MUX2_X1 _26483_ (.A(_08275_),
    .B(\cs_registers_i.mscratch_q[11] ),
    .S(_08743_),
    .Z(_01982_));
 MUX2_X1 _26484_ (.A(_08444_),
    .B(\cs_registers_i.mscratch_q[12] ),
    .S(_08743_),
    .Z(_01983_));
 MUX2_X1 _26485_ (.A(_07569_),
    .B(\cs_registers_i.mscratch_q[13] ),
    .S(_08743_),
    .Z(_01984_));
 MUX2_X1 _26486_ (.A(_07579_),
    .B(\cs_registers_i.mscratch_q[14] ),
    .S(_08743_),
    .Z(_01985_));
 MUX2_X1 _26487_ (.A(_08299_),
    .B(\cs_registers_i.mscratch_q[15] ),
    .S(_08743_),
    .Z(_01986_));
 MUX2_X1 _26488_ (.A(_07600_),
    .B(\cs_registers_i.mscratch_q[16] ),
    .S(_08743_),
    .Z(_01987_));
 NAND2_X1 _26489_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(_08744_),
    .ZN(_08747_));
 OAI21_X1 _26490_ (.A(_08747_),
    .B1(_08746_),
    .B2(_08312_),
    .ZN(_01988_));
 MUX2_X1 _26491_ (.A(_07914_),
    .B(\cs_registers_i.mscratch_q[18] ),
    .S(_08743_),
    .Z(_01989_));
 NAND2_X1 _26492_ (.A1(\cs_registers_i.mscratch_q[19] ),
    .A2(_08744_),
    .ZN(_08748_));
 OAI21_X1 _26493_ (.A(_08748_),
    .B1(_08746_),
    .B2(_07624_),
    .ZN(_01990_));
 NAND2_X1 _26494_ (.A1(\cs_registers_i.mscratch_q[1] ),
    .A2(_08744_),
    .ZN(_08749_));
 OAI21_X1 _26495_ (.A(_08749_),
    .B1(_08746_),
    .B2(_07635_),
    .ZN(_01991_));
 NAND2_X1 _26496_ (.A1(\cs_registers_i.mscratch_q[20] ),
    .A2(_08744_),
    .ZN(_08750_));
 OAI21_X1 _26497_ (.A(_08750_),
    .B1(_08746_),
    .B2(_07640_),
    .ZN(_01992_));
 MUX2_X1 _26498_ (.A(_08343_),
    .B(\cs_registers_i.mscratch_q[21] ),
    .S(_08743_),
    .Z(_01993_));
 NAND2_X1 _26499_ (.A1(\cs_registers_i.mscratch_q[22] ),
    .A2(_08744_),
    .ZN(_08751_));
 OAI21_X1 _26500_ (.A(_08751_),
    .B1(_08746_),
    .B2(_07657_),
    .ZN(_01994_));
 MUX2_X1 _26501_ (.A(_08355_),
    .B(\cs_registers_i.mscratch_q[23] ),
    .S(_08743_),
    .Z(_01995_));
 BUF_X4 _26502_ (.A(_08742_),
    .Z(_08752_));
 MUX2_X1 _26503_ (.A(_08149_),
    .B(\cs_registers_i.mscratch_q[24] ),
    .S(_08752_),
    .Z(_01996_));
 MUX2_X1 _26504_ (.A(_07689_),
    .B(\cs_registers_i.mscratch_q[25] ),
    .S(_08752_),
    .Z(_01997_));
 NAND2_X1 _26505_ (.A1(\cs_registers_i.mscratch_q[26] ),
    .A2(_08744_),
    .ZN(_08753_));
 OAI21_X1 _26506_ (.A(_08753_),
    .B1(_08746_),
    .B2(_08163_),
    .ZN(_01998_));
 NAND2_X1 _26507_ (.A1(\cs_registers_i.mscratch_q[27] ),
    .A2(_08744_),
    .ZN(_08754_));
 OAI21_X1 _26508_ (.A(_08754_),
    .B1(_08746_),
    .B2(_07709_),
    .ZN(_01999_));
 MUX2_X1 _26509_ (.A(_07718_),
    .B(\cs_registers_i.mscratch_q[28] ),
    .S(_08752_),
    .Z(_02000_));
 NAND2_X1 _26510_ (.A1(\cs_registers_i.mscratch_q[29] ),
    .A2(_08744_),
    .ZN(_08755_));
 OAI21_X1 _26511_ (.A(_08755_),
    .B1(_08746_),
    .B2(_07728_),
    .ZN(_02001_));
 MUX2_X1 _26512_ (.A(_07493_),
    .B(\cs_registers_i.mscratch_q[2] ),
    .S(_08752_),
    .Z(_02002_));
 NAND2_X1 _26513_ (.A1(\cs_registers_i.mscratch_q[30] ),
    .A2(_08744_),
    .ZN(_08756_));
 OAI21_X1 _26514_ (.A(_08756_),
    .B1(_08746_),
    .B2(_07983_),
    .ZN(_02003_));
 MUX2_X1 _26515_ (.A(_08405_),
    .B(\cs_registers_i.mscratch_q[31] ),
    .S(_08752_),
    .Z(_02004_));
 MUX2_X1 _26516_ (.A(_08224_),
    .B(\cs_registers_i.mscratch_q[3] ),
    .S(_08752_),
    .Z(_02005_));
 MUX2_X1 _26517_ (.A(_08231_),
    .B(\cs_registers_i.mscratch_q[4] ),
    .S(_08752_),
    .Z(_02006_));
 MUX2_X1 _26518_ (.A(_07810_),
    .B(\cs_registers_i.mscratch_q[5] ),
    .S(_08752_),
    .Z(_02007_));
 MUX2_X1 _26519_ (.A(_08243_),
    .B(\cs_registers_i.mscratch_q[6] ),
    .S(_08752_),
    .Z(_02008_));
 MUX2_X1 _26520_ (.A(_08250_),
    .B(\cs_registers_i.mscratch_q[7] ),
    .S(_08752_),
    .Z(_02009_));
 MUX2_X1 _26521_ (.A(_07844_),
    .B(\cs_registers_i.mscratch_q[8] ),
    .S(_08742_),
    .Z(_02010_));
 MUX2_X1 _26522_ (.A(_07854_),
    .B(\cs_registers_i.mscratch_q[9] ),
    .S(_08742_),
    .Z(_02011_));
 CLKBUF_X3 _26523_ (.A(_08596_),
    .Z(_08757_));
 MUX2_X1 _26524_ (.A(\cs_registers_i.mcause_q[0] ),
    .B(\cs_registers_i.mstack_cause_q[0] ),
    .S(_08757_),
    .Z(_02012_));
 MUX2_X1 _26525_ (.A(\cs_registers_i.mcause_q[1] ),
    .B(\cs_registers_i.mstack_cause_q[1] ),
    .S(_08757_),
    .Z(_02013_));
 MUX2_X1 _26526_ (.A(\cs_registers_i.mcause_q[2] ),
    .B(\cs_registers_i.mstack_cause_q[2] ),
    .S(_08757_),
    .Z(_02014_));
 MUX2_X1 _26527_ (.A(\cs_registers_i.mcause_q[3] ),
    .B(\cs_registers_i.mstack_cause_q[3] ),
    .S(_08757_),
    .Z(_02015_));
 MUX2_X1 _26528_ (.A(\cs_registers_i.mcause_q[4] ),
    .B(\cs_registers_i.mstack_cause_q[4] ),
    .S(_08757_),
    .Z(_02016_));
 MUX2_X1 _26529_ (.A(\cs_registers_i.mcause_q[5] ),
    .B(\cs_registers_i.mstack_cause_q[5] ),
    .S(_08757_),
    .Z(_02017_));
 MUX2_X1 _26530_ (.A(\cs_registers_i.mstack_d[0] ),
    .B(\cs_registers_i.mstack_q[0] ),
    .S(_08757_),
    .Z(_02018_));
 MUX2_X1 _26531_ (.A(\cs_registers_i.mstack_d[1] ),
    .B(\cs_registers_i.mstack_q[1] ),
    .S(_08757_),
    .Z(_02019_));
 BUF_X4 _26532_ (.A(_08596_),
    .Z(_08758_));
 MUX2_X1 _26533_ (.A(\cs_registers_i.mstack_d[2] ),
    .B(\cs_registers_i.mstack_q[2] ),
    .S(_08758_),
    .Z(_02020_));
 MUX2_X1 _26534_ (.A(\cs_registers_i.csr_mepc_o[0] ),
    .B(\cs_registers_i.mstack_epc_q[0] ),
    .S(_08758_),
    .Z(_02021_));
 MUX2_X1 _26535_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(\cs_registers_i.mstack_epc_q[10] ),
    .S(_08758_),
    .Z(_02022_));
 MUX2_X1 _26536_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(\cs_registers_i.mstack_epc_q[11] ),
    .S(_08758_),
    .Z(_02023_));
 MUX2_X1 _26537_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(\cs_registers_i.mstack_epc_q[12] ),
    .S(_08758_),
    .Z(_02024_));
 MUX2_X1 _26538_ (.A(\cs_registers_i.csr_mepc_o[13] ),
    .B(\cs_registers_i.mstack_epc_q[13] ),
    .S(_08758_),
    .Z(_02025_));
 MUX2_X1 _26539_ (.A(\cs_registers_i.csr_mepc_o[14] ),
    .B(\cs_registers_i.mstack_epc_q[14] ),
    .S(_08758_),
    .Z(_02026_));
 MUX2_X1 _26540_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(\cs_registers_i.mstack_epc_q[15] ),
    .S(_08758_),
    .Z(_02027_));
 MUX2_X1 _26541_ (.A(\cs_registers_i.csr_mepc_o[16] ),
    .B(\cs_registers_i.mstack_epc_q[16] ),
    .S(_08758_),
    .Z(_02028_));
 MUX2_X1 _26542_ (.A(\cs_registers_i.csr_mepc_o[17] ),
    .B(\cs_registers_i.mstack_epc_q[17] ),
    .S(_08758_),
    .Z(_02029_));
 BUF_X4 _26543_ (.A(_08595_),
    .Z(_08759_));
 MUX2_X1 _26544_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(\cs_registers_i.mstack_epc_q[18] ),
    .S(_08759_),
    .Z(_02030_));
 MUX2_X1 _26545_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(\cs_registers_i.mstack_epc_q[19] ),
    .S(_08759_),
    .Z(_02031_));
 MUX2_X1 _26546_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(\cs_registers_i.mstack_epc_q[1] ),
    .S(_08759_),
    .Z(_02032_));
 MUX2_X1 _26547_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(\cs_registers_i.mstack_epc_q[20] ),
    .S(_08759_),
    .Z(_02033_));
 MUX2_X1 _26548_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(\cs_registers_i.mstack_epc_q[21] ),
    .S(_08759_),
    .Z(_02034_));
 MUX2_X1 _26549_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(\cs_registers_i.mstack_epc_q[22] ),
    .S(_08759_),
    .Z(_02035_));
 MUX2_X1 _26550_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(\cs_registers_i.mstack_epc_q[23] ),
    .S(_08759_),
    .Z(_02036_));
 MUX2_X1 _26551_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(\cs_registers_i.mstack_epc_q[24] ),
    .S(_08759_),
    .Z(_02037_));
 MUX2_X1 _26552_ (.A(\cs_registers_i.csr_mepc_o[25] ),
    .B(\cs_registers_i.mstack_epc_q[25] ),
    .S(_08759_),
    .Z(_02038_));
 MUX2_X1 _26553_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(\cs_registers_i.mstack_epc_q[26] ),
    .S(_08759_),
    .Z(_02039_));
 BUF_X4 _26554_ (.A(_08595_),
    .Z(_08760_));
 MUX2_X1 _26555_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(\cs_registers_i.mstack_epc_q[27] ),
    .S(_08760_),
    .Z(_02040_));
 MUX2_X1 _26556_ (.A(\cs_registers_i.csr_mepc_o[28] ),
    .B(\cs_registers_i.mstack_epc_q[28] ),
    .S(_08760_),
    .Z(_02041_));
 MUX2_X1 _26557_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(\cs_registers_i.mstack_epc_q[29] ),
    .S(_08760_),
    .Z(_02042_));
 MUX2_X1 _26558_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .B(\cs_registers_i.mstack_epc_q[2] ),
    .S(_08760_),
    .Z(_02043_));
 MUX2_X1 _26559_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(\cs_registers_i.mstack_epc_q[30] ),
    .S(_08760_),
    .Z(_02044_));
 MUX2_X1 _26560_ (.A(\cs_registers_i.csr_mepc_o[31] ),
    .B(\cs_registers_i.mstack_epc_q[31] ),
    .S(_08760_),
    .Z(_02045_));
 MUX2_X1 _26561_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(\cs_registers_i.mstack_epc_q[3] ),
    .S(_08760_),
    .Z(_02046_));
 MUX2_X1 _26562_ (.A(\cs_registers_i.csr_mepc_o[4] ),
    .B(\cs_registers_i.mstack_epc_q[4] ),
    .S(_08760_),
    .Z(_02047_));
 MUX2_X1 _26563_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .B(\cs_registers_i.mstack_epc_q[5] ),
    .S(_08760_),
    .Z(_02048_));
 MUX2_X1 _26564_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(\cs_registers_i.mstack_epc_q[6] ),
    .S(_08760_),
    .Z(_02049_));
 MUX2_X1 _26565_ (.A(\cs_registers_i.csr_mepc_o[7] ),
    .B(\cs_registers_i.mstack_epc_q[7] ),
    .S(_08596_),
    .Z(_02050_));
 MUX2_X1 _26566_ (.A(\cs_registers_i.csr_mepc_o[8] ),
    .B(\cs_registers_i.mstack_epc_q[8] ),
    .S(_08596_),
    .Z(_02051_));
 MUX2_X1 _26567_ (.A(\cs_registers_i.csr_mepc_o[9] ),
    .B(\cs_registers_i.mstack_epc_q[9] ),
    .S(_08596_),
    .Z(_02052_));
 NAND2_X2 _26568_ (.A1(_05487_),
    .A2(_07489_),
    .ZN(_08761_));
 MUX2_X1 _26569_ (.A(_08343_),
    .B(\cs_registers_i.csr_mstatus_tw_o ),
    .S(_08761_),
    .Z(_02053_));
 NAND2_X1 _26570_ (.A1(\cs_registers_i.mstatus_q[1] ),
    .A2(_08761_),
    .ZN(_08762_));
 OAI21_X1 _26571_ (.A(_08762_),
    .B1(_08761_),
    .B2(_08312_),
    .ZN(_02054_));
 NOR2_X2 _26572_ (.A1(_03954_),
    .A2(_08615_),
    .ZN(_08763_));
 NOR2_X1 _26573_ (.A1(_06797_),
    .A2(_08763_),
    .ZN(_08764_));
 NAND3_X1 _26574_ (.A1(_03487_),
    .A2(_04261_),
    .A3(_05487_),
    .ZN(_08765_));
 NAND2_X1 _26575_ (.A1(_08764_),
    .A2(_08765_),
    .ZN(_08766_));
 AOI22_X1 _26576_ (.A1(\cs_registers_i.mstack_q[0] ),
    .A2(_08588_),
    .B1(_08633_),
    .B2(_03462_),
    .ZN(_08767_));
 INV_X1 _26577_ (.A(_08767_),
    .ZN(_08768_));
 AOI21_X1 _26578_ (.A(_08761_),
    .B1(_07554_),
    .B2(_07535_),
    .ZN(_08769_));
 OAI21_X1 _26579_ (.A(_08766_),
    .B1(_08768_),
    .B2(_08769_),
    .ZN(_08770_));
 AOI21_X1 _26580_ (.A(_06797_),
    .B1(_08763_),
    .B2(_08633_),
    .ZN(_08771_));
 NAND2_X1 _26581_ (.A1(_08761_),
    .A2(_08771_),
    .ZN(_08772_));
 INV_X1 _26582_ (.A(\cs_registers_i.mstack_d[0] ),
    .ZN(_08773_));
 OAI21_X1 _26583_ (.A(_08770_),
    .B1(_08772_),
    .B2(_08773_),
    .ZN(_02055_));
 BUF_X4 _26584_ (.A(_08620_),
    .Z(_08774_));
 AOI22_X1 _26585_ (.A1(\cs_registers_i.mstack_q[1] ),
    .A2(_08588_),
    .B1(_08774_),
    .B2(_03463_),
    .ZN(_08775_));
 INV_X1 _26586_ (.A(_08775_),
    .ZN(_08776_));
 OAI21_X1 _26587_ (.A(_08766_),
    .B1(_08769_),
    .B2(_08776_),
    .ZN(_08777_));
 INV_X1 _26588_ (.A(\cs_registers_i.mstack_d[1] ),
    .ZN(_08778_));
 OAI21_X1 _26589_ (.A(_08777_),
    .B1(_08772_),
    .B2(_08778_),
    .ZN(_02056_));
 INV_X1 _26590_ (.A(\cs_registers_i.mstack_q[2] ),
    .ZN(_08779_));
 NAND3_X1 _26591_ (.A1(_03870_),
    .A2(_08779_),
    .A3(_06803_),
    .ZN(_08780_));
 AOI22_X1 _26592_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_08633_),
    .B1(_08780_),
    .B2(_06797_),
    .ZN(_08781_));
 OAI21_X1 _26593_ (.A(_08781_),
    .B1(_08761_),
    .B2(_07828_),
    .ZN(_08782_));
 NAND2_X1 _26594_ (.A1(_08766_),
    .A2(_08782_),
    .ZN(_08783_));
 AOI21_X1 _26595_ (.A(_08633_),
    .B1(_08588_),
    .B2(_08779_),
    .ZN(_08784_));
 AOI22_X1 _26596_ (.A1(_08764_),
    .A2(_08765_),
    .B1(_08784_),
    .B2(_08761_),
    .ZN(_08785_));
 INV_X1 _26597_ (.A(\cs_registers_i.mstack_d[2] ),
    .ZN(_08786_));
 OAI21_X1 _26598_ (.A(_08783_),
    .B1(_08785_),
    .B2(_08786_),
    .ZN(_02057_));
 NOR2_X1 _26599_ (.A1(_07791_),
    .A2(_08761_),
    .ZN(_08787_));
 AOI21_X1 _26600_ (.A(_08787_),
    .B1(_06797_),
    .B2(\cs_registers_i.mstack_d[2] ),
    .ZN(_08788_));
 INV_X1 _26601_ (.A(\cs_registers_i.csr_mstatus_mie_o ),
    .ZN(_08789_));
 OAI21_X1 _26602_ (.A(_08788_),
    .B1(_08766_),
    .B2(_08789_),
    .ZN(_02058_));
 AND4_X1 _26603_ (.A1(_08600_),
    .A2(_03842_),
    .A3(_03610_),
    .A4(_03837_),
    .ZN(_08790_));
 BUF_X4 _26604_ (.A(_08790_),
    .Z(_08791_));
 BUF_X4 _26605_ (.A(_08791_),
    .Z(_08792_));
 MUX2_X2 _26606_ (.A(_10291_),
    .B(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(_10338_),
    .Z(_08793_));
 AOI22_X1 _26607_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(_08792_),
    .B1(_08793_),
    .B2(_08604_),
    .ZN(_08794_));
 OR3_X1 _26608_ (.A1(_08595_),
    .A2(_08634_),
    .A3(_08794_),
    .ZN(_08795_));
 CLKBUF_X3 _26609_ (.A(_08647_),
    .Z(_08796_));
 OAI21_X1 _26610_ (.A(_08795_),
    .B1(_08796_),
    .B2(_07482_),
    .ZN(_08797_));
 AOI21_X4 _26611_ (.A(_08763_),
    .B1(_07488_),
    .B2(_04521_),
    .ZN(_08798_));
 BUF_X4 _26612_ (.A(_08798_),
    .Z(_08799_));
 MUX2_X1 _26613_ (.A(_08797_),
    .B(\cs_registers_i.mtval_q[0] ),
    .S(_08799_),
    .Z(_02059_));
 CLKBUF_X3 _26614_ (.A(_06989_),
    .Z(_08800_));
 BUF_X4 _26615_ (.A(_03607_),
    .Z(_08801_));
 CLKBUF_X3 _26616_ (.A(_08801_),
    .Z(_08802_));
 BUF_X4 _26617_ (.A(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_08803_));
 NAND3_X1 _26618_ (.A1(_10675_),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(_08803_),
    .ZN(_08804_));
 NAND3_X1 _26619_ (.A1(_11517_),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(\cs_registers_i.pc_id_i[5] ),
    .ZN(_08805_));
 NOR2_X1 _26620_ (.A1(_11673_),
    .A2(_08805_),
    .ZN(_08806_));
 NAND2_X1 _26621_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_08806_),
    .ZN(_08807_));
 NOR2_X2 _26622_ (.A1(_08804_),
    .A2(_08807_),
    .ZN(_08808_));
 NAND3_X1 _26623_ (.A1(_11788_),
    .A2(_11826_),
    .A3(_08808_),
    .ZN(_08809_));
 XNOR2_X1 _26624_ (.A(_00038_),
    .B(_08809_),
    .ZN(_08810_));
 NAND2_X1 _26625_ (.A1(_08802_),
    .A2(_08810_),
    .ZN(_08811_));
 INV_X1 _26626_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .ZN(_08812_));
 BUF_X4 _26627_ (.A(_10338_),
    .Z(_08813_));
 MUX2_X2 _26628_ (.A(_00036_),
    .B(_00037_),
    .S(_08813_),
    .Z(_08814_));
 BUF_X4 _26629_ (.A(_08601_),
    .Z(_08815_));
 OAI221_X2 _26630_ (.A(_08599_),
    .B1(_08603_),
    .B2(_08812_),
    .C1(_08814_),
    .C2(_08815_),
    .ZN(_08816_));
 NAND4_X2 _26631_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08811_),
    .A4(_08816_),
    .ZN(_08817_));
 OAI21_X1 _26632_ (.A(_08817_),
    .B1(_08796_),
    .B2(_07525_),
    .ZN(_08818_));
 MUX2_X1 _26633_ (.A(_08818_),
    .B(\cs_registers_i.mtval_q[10] ),
    .S(_08799_),
    .Z(_02060_));
 CLKBUF_X3 _26634_ (.A(_08620_),
    .Z(_08819_));
 NAND2_X1 _26635_ (.A1(_08803_),
    .A2(_15536_),
    .ZN(_08820_));
 NOR2_X2 _26636_ (.A1(_08807_),
    .A2(_08820_),
    .ZN(_08821_));
 NAND4_X1 _26637_ (.A1(_11788_),
    .A2(_11826_),
    .A3(\cs_registers_i.pc_id_i[10] ),
    .A4(_08821_),
    .ZN(_08822_));
 XNOR2_X1 _26638_ (.A(_00041_),
    .B(_08822_),
    .ZN(_08823_));
 NAND2_X1 _26639_ (.A1(_08802_),
    .A2(_08823_),
    .ZN(_08824_));
 INV_X1 _26640_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .ZN(_08825_));
 MUX2_X2 _26641_ (.A(_04603_),
    .B(_00040_),
    .S(_08813_),
    .Z(_08826_));
 OAI221_X2 _26642_ (.A(_08599_),
    .B1(_08603_),
    .B2(_08825_),
    .C1(_08826_),
    .C2(_08815_),
    .ZN(_08827_));
 NAND4_X2 _26643_ (.A1(_08800_),
    .A2(_08819_),
    .A3(_08824_),
    .A4(_08827_),
    .ZN(_08828_));
 OAI21_X1 _26644_ (.A(_08828_),
    .B1(_08796_),
    .B2(_07535_),
    .ZN(_08829_));
 MUX2_X1 _26645_ (.A(_08829_),
    .B(\cs_registers_i.mtval_q[11] ),
    .S(_08799_),
    .Z(_02061_));
 AND4_X2 _26646_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_11788_),
    .A3(_11826_),
    .A4(\cs_registers_i.pc_id_i[10] ),
    .ZN(_08830_));
 NAND2_X1 _26647_ (.A1(_08808_),
    .A2(_08830_),
    .ZN(_08831_));
 XNOR2_X1 _26648_ (.A(_00043_),
    .B(_08831_),
    .ZN(_08832_));
 NAND2_X1 _26649_ (.A1(_08802_),
    .A2(_08832_),
    .ZN(_08833_));
 INV_X1 _26650_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .ZN(_08834_));
 MUX2_X2 _26651_ (.A(_00176_),
    .B(_00042_),
    .S(_08813_),
    .Z(_08835_));
 OAI221_X2 _26652_ (.A(_08599_),
    .B1(_08603_),
    .B2(_08834_),
    .C1(_08835_),
    .C2(_08815_),
    .ZN(_08836_));
 NAND4_X2 _26653_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08833_),
    .A4(_08836_),
    .ZN(_08837_));
 OAI21_X1 _26654_ (.A(_08837_),
    .B1(_08796_),
    .B2(_07554_),
    .ZN(_08838_));
 CLKBUF_X3 _26655_ (.A(_08798_),
    .Z(_08839_));
 MUX2_X1 _26656_ (.A(_08838_),
    .B(\cs_registers_i.mtval_q[12] ),
    .S(_08839_),
    .Z(_02062_));
 NAND2_X1 _26657_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(_08799_),
    .ZN(_08840_));
 INV_X1 _26658_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .ZN(_08841_));
 MUX2_X2 _26659_ (.A(_00175_),
    .B(_00044_),
    .S(_10338_),
    .Z(_08842_));
 OAI221_X2 _26660_ (.A(_08598_),
    .B1(_08602_),
    .B2(_08841_),
    .C1(_08842_),
    .C2(_08601_),
    .ZN(_08843_));
 NAND3_X4 _26661_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_08821_),
    .A3(_08830_),
    .ZN(_08844_));
 XOR2_X2 _26662_ (.A(_00045_),
    .B(_08844_),
    .Z(_08845_));
 OAI21_X1 _26663_ (.A(_08843_),
    .B1(_08845_),
    .B2(_08599_),
    .ZN(_08846_));
 NOR3_X1 _26664_ (.A1(_08621_),
    .A2(_08596_),
    .A3(_08846_),
    .ZN(_08847_));
 AOI21_X1 _26665_ (.A(_08847_),
    .B1(_08757_),
    .B2(_07569_),
    .ZN(_08848_));
 OAI21_X1 _26666_ (.A(_08840_),
    .B1(_08848_),
    .B2(_08799_),
    .ZN(_02063_));
 NAND3_X2 _26667_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_08808_),
    .A3(_08830_),
    .ZN(_08849_));
 INV_X1 _26668_ (.A(_08849_),
    .ZN(_08850_));
 NAND2_X1 _26669_ (.A1(_12076_),
    .A2(_08850_),
    .ZN(_08851_));
 XNOR2_X1 _26670_ (.A(_00047_),
    .B(_08851_),
    .ZN(_08852_));
 NAND2_X1 _26671_ (.A1(_08802_),
    .A2(_08852_),
    .ZN(_08853_));
 BUF_X4 _26672_ (.A(_08598_),
    .Z(_08854_));
 INV_X1 _26673_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .ZN(_08855_));
 MUX2_X2 _26674_ (.A(_10522_),
    .B(_00046_),
    .S(_08813_),
    .Z(_08856_));
 OAI221_X2 _26675_ (.A(_08854_),
    .B1(_08603_),
    .B2(_08855_),
    .C1(_08856_),
    .C2(_08815_),
    .ZN(_08857_));
 NAND4_X2 _26676_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08853_),
    .A4(_08857_),
    .ZN(_08858_));
 OAI21_X1 _26677_ (.A(_08858_),
    .B1(_08796_),
    .B2(_08089_),
    .ZN(_08859_));
 MUX2_X1 _26678_ (.A(_08859_),
    .B(\cs_registers_i.mtval_q[14] ),
    .S(_08839_),
    .Z(_02064_));
 INV_X1 _26679_ (.A(_08844_),
    .ZN(_08860_));
 NAND3_X1 _26680_ (.A1(_12076_),
    .A2(_12179_),
    .A3(_08860_),
    .ZN(_08861_));
 XNOR2_X1 _26681_ (.A(_00049_),
    .B(_08861_),
    .ZN(_08862_));
 NAND2_X1 _26682_ (.A1(_08802_),
    .A2(_08862_),
    .ZN(_08863_));
 INV_X1 _26683_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .ZN(_08864_));
 MUX2_X1 _26684_ (.A(_00184_),
    .B(_00048_),
    .S(_08813_),
    .Z(_08865_));
 OAI221_X2 _26685_ (.A(_08854_),
    .B1(_08603_),
    .B2(_08864_),
    .C1(_08865_),
    .C2(_08815_),
    .ZN(_08866_));
 NAND4_X2 _26686_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08863_),
    .A4(_08866_),
    .ZN(_08867_));
 OAI21_X1 _26687_ (.A(_08867_),
    .B1(_08796_),
    .B2(_07585_),
    .ZN(_08868_));
 MUX2_X1 _26688_ (.A(_08868_),
    .B(\cs_registers_i.mtval_q[15] ),
    .S(_08839_),
    .Z(_02065_));
 NOR2_X4 _26689_ (.A1(_10338_),
    .A2(_03842_),
    .ZN(_08869_));
 BUF_X4 _26690_ (.A(_08869_),
    .Z(_08870_));
 AOI221_X2 _26691_ (.A(_08801_),
    .B1(_08792_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .C1(_08870_),
    .C2(_10759_),
    .ZN(_08871_));
 NAND3_X1 _26692_ (.A1(_12076_),
    .A2(_12179_),
    .A3(\cs_registers_i.pc_id_i[15] ),
    .ZN(_08872_));
 NOR2_X1 _26693_ (.A1(_08849_),
    .A2(_08872_),
    .ZN(_08873_));
 XOR2_X2 _26694_ (.A(_00050_),
    .B(_08873_),
    .Z(_08874_));
 BUF_X4 _26695_ (.A(_08801_),
    .Z(_08875_));
 AOI21_X2 _26696_ (.A(_08871_),
    .B1(_08874_),
    .B2(_08875_),
    .ZN(_08876_));
 NAND3_X2 _26697_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08876_),
    .ZN(_08877_));
 OAI21_X1 _26698_ (.A(_08877_),
    .B1(_08796_),
    .B2(_08100_),
    .ZN(_08878_));
 MUX2_X1 _26699_ (.A(_08878_),
    .B(\cs_registers_i.mtval_q[16] ),
    .S(_08839_),
    .Z(_02066_));
 AOI221_X2 _26700_ (.A(_08801_),
    .B1(_08792_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .C1(_08870_),
    .C2(_10752_),
    .ZN(_08879_));
 NOR2_X2 _26701_ (.A1(_12352_),
    .A2(_08872_),
    .ZN(_08880_));
 NAND2_X1 _26702_ (.A1(_08860_),
    .A2(_08880_),
    .ZN(_08881_));
 XNOR2_X1 _26703_ (.A(_00051_),
    .B(_08881_),
    .ZN(_08882_));
 AOI21_X1 _26704_ (.A(_08879_),
    .B1(_08882_),
    .B2(_08875_),
    .ZN(_08883_));
 NAND3_X1 _26705_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08883_),
    .ZN(_08884_));
 OAI21_X1 _26706_ (.A(_08884_),
    .B1(_08796_),
    .B2(_08312_),
    .ZN(_08885_));
 MUX2_X1 _26707_ (.A(_08885_),
    .B(\cs_registers_i.mtval_q[17] ),
    .S(_08839_),
    .Z(_02067_));
 AOI221_X2 _26708_ (.A(_08801_),
    .B1(_08792_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .C1(_08870_),
    .C2(_10767_),
    .ZN(_08886_));
 NAND3_X1 _26709_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_08850_),
    .A3(_08880_),
    .ZN(_08887_));
 XNOR2_X1 _26710_ (.A(_00052_),
    .B(_08887_),
    .ZN(_08888_));
 AOI21_X1 _26711_ (.A(_08886_),
    .B1(_08888_),
    .B2(_08875_),
    .ZN(_08889_));
 NAND3_X1 _26712_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08889_),
    .ZN(_08890_));
 OAI21_X1 _26713_ (.A(_08890_),
    .B1(_08796_),
    .B2(_07616_),
    .ZN(_08891_));
 MUX2_X1 _26714_ (.A(_08891_),
    .B(\cs_registers_i.mtval_q[18] ),
    .S(_08839_),
    .Z(_02068_));
 AOI221_X1 _26715_ (.A(_08801_),
    .B1(_08792_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .C1(_08870_),
    .C2(_10750_),
    .ZN(_08892_));
 NAND3_X4 _26716_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(\cs_registers_i.pc_id_i[18] ),
    .A3(_08880_),
    .ZN(_08893_));
 NOR2_X1 _26717_ (.A1(_08844_),
    .A2(_08893_),
    .ZN(_08894_));
 XOR2_X1 _26718_ (.A(_00053_),
    .B(_08894_),
    .Z(_08895_));
 AOI21_X1 _26719_ (.A(_08892_),
    .B1(_08895_),
    .B2(_08875_),
    .ZN(_08896_));
 NAND3_X1 _26720_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08896_),
    .ZN(_08897_));
 OAI21_X1 _26721_ (.A(_08897_),
    .B1(_08796_),
    .B2(_07624_),
    .ZN(_08898_));
 MUX2_X1 _26722_ (.A(_08898_),
    .B(\cs_registers_i.mtval_q[19] ),
    .S(_08839_),
    .Z(_02069_));
 INV_X1 _26723_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .ZN(_08899_));
 MUX2_X2 _26724_ (.A(_00013_),
    .B(_00014_),
    .S(_08813_),
    .Z(_08900_));
 OAI221_X1 _26725_ (.A(_08599_),
    .B1(_08603_),
    .B2(_08899_),
    .C1(_08900_),
    .C2(_08815_),
    .ZN(_08901_));
 XNOR2_X1 _26726_ (.A(_10675_),
    .B(_08803_),
    .ZN(_08902_));
 NAND2_X1 _26727_ (.A1(_08802_),
    .A2(_08902_),
    .ZN(_08903_));
 NAND4_X1 _26728_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08901_),
    .A4(_08903_),
    .ZN(_08904_));
 CLKBUF_X3 _26729_ (.A(_08647_),
    .Z(_08905_));
 OAI21_X1 _26730_ (.A(_08904_),
    .B1(_08905_),
    .B2(_07635_),
    .ZN(_08906_));
 MUX2_X1 _26731_ (.A(_08906_),
    .B(\cs_registers_i.mtval_q[1] ),
    .S(_08839_),
    .Z(_02070_));
 AOI221_X2 _26732_ (.A(_08801_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .C1(_08870_),
    .C2(_11935_),
    .ZN(_08907_));
 NOR2_X1 _26733_ (.A1(_08849_),
    .A2(_08893_),
    .ZN(_08908_));
 NAND2_X1 _26734_ (.A1(_12590_),
    .A2(_08908_),
    .ZN(_08909_));
 XNOR2_X1 _26735_ (.A(_00054_),
    .B(_08909_),
    .ZN(_08910_));
 AOI21_X1 _26736_ (.A(_08907_),
    .B1(_08910_),
    .B2(_08875_),
    .ZN(_08911_));
 NAND3_X1 _26737_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08911_),
    .ZN(_08912_));
 OAI21_X1 _26738_ (.A(_08912_),
    .B1(_08905_),
    .B2(_07640_),
    .ZN(_08913_));
 MUX2_X1 _26739_ (.A(_08913_),
    .B(\cs_registers_i.mtval_q[20] ),
    .S(_08839_),
    .Z(_02071_));
 AOI221_X2 _26740_ (.A(_08801_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .C1(_08869_),
    .C2(_12034_),
    .ZN(_08914_));
 NAND3_X1 _26741_ (.A1(_12590_),
    .A2(_12685_),
    .A3(_08894_),
    .ZN(_08915_));
 XNOR2_X1 _26742_ (.A(_00055_),
    .B(_08915_),
    .ZN(_08916_));
 AOI21_X1 _26743_ (.A(_08914_),
    .B1(_08916_),
    .B2(_08875_),
    .ZN(_08917_));
 NAND3_X1 _26744_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08917_),
    .ZN(_08918_));
 OAI21_X1 _26745_ (.A(_08918_),
    .B1(_08905_),
    .B2(_07651_),
    .ZN(_08919_));
 MUX2_X1 _26746_ (.A(_08919_),
    .B(\cs_registers_i.mtval_q[21] ),
    .S(_08839_),
    .Z(_02072_));
 AOI221_X2 _26747_ (.A(_03607_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .C1(_08869_),
    .C2(_11989_),
    .ZN(_08920_));
 NAND4_X1 _26748_ (.A1(_12590_),
    .A2(_12685_),
    .A3(\cs_registers_i.pc_id_i[21] ),
    .A4(_08908_),
    .ZN(_08921_));
 XNOR2_X1 _26749_ (.A(_00056_),
    .B(_08921_),
    .ZN(_08922_));
 AOI21_X1 _26750_ (.A(_08920_),
    .B1(_08922_),
    .B2(_08875_),
    .ZN(_08923_));
 NAND3_X1 _26751_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08923_),
    .ZN(_08924_));
 OAI21_X2 _26752_ (.A(_08924_),
    .B1(_08905_),
    .B2(_07657_),
    .ZN(_08925_));
 BUF_X4 _26753_ (.A(_08798_),
    .Z(_08926_));
 MUX2_X1 _26754_ (.A(_08925_),
    .B(\cs_registers_i.mtval_q[22] ),
    .S(_08926_),
    .Z(_02073_));
 AOI221_X2 _26755_ (.A(_03607_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .C1(_08869_),
    .C2(_12041_),
    .ZN(_08927_));
 NAND4_X4 _26756_ (.A1(_12590_),
    .A2(_12685_),
    .A3(\cs_registers_i.pc_id_i[21] ),
    .A4(\cs_registers_i.pc_id_i[22] ),
    .ZN(_08928_));
 NOR3_X4 _26757_ (.A1(_08844_),
    .A2(_08893_),
    .A3(_08928_),
    .ZN(_08929_));
 XOR2_X1 _26758_ (.A(_00057_),
    .B(_08929_),
    .Z(_08930_));
 AOI21_X1 _26759_ (.A(_08927_),
    .B1(_08930_),
    .B2(_08875_),
    .ZN(_08931_));
 NAND3_X1 _26760_ (.A1(_08800_),
    .A2(_08774_),
    .A3(_08931_),
    .ZN(_08932_));
 OAI21_X1 _26761_ (.A(_08932_),
    .B1(_08905_),
    .B2(_07669_),
    .ZN(_08933_));
 MUX2_X1 _26762_ (.A(_08933_),
    .B(\cs_registers_i.mtval_q[23] ),
    .S(_08926_),
    .Z(_02074_));
 AOI221_X2 _26763_ (.A(_03607_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .C1(_08869_),
    .C2(_11929_),
    .ZN(_08934_));
 NOR3_X2 _26764_ (.A1(_08849_),
    .A2(_08893_),
    .A3(_08928_),
    .ZN(_08935_));
 NAND2_X1 _26765_ (.A1(_12935_),
    .A2(_08935_),
    .ZN(_08936_));
 XNOR2_X1 _26766_ (.A(_00058_),
    .B(_08936_),
    .ZN(_08937_));
 AOI21_X2 _26767_ (.A(_08934_),
    .B1(_08937_),
    .B2(_08875_),
    .ZN(_08938_));
 NOR2_X2 _26768_ (.A1(_08621_),
    .A2(_08592_),
    .ZN(_08939_));
 AOI221_X2 _26769_ (.A(_08798_),
    .B1(_08938_),
    .B2(_08939_),
    .C1(_08595_),
    .C2(_08149_),
    .ZN(_08940_));
 INV_X1 _26770_ (.A(\cs_registers_i.mtval_q[24] ),
    .ZN(_08941_));
 AOI21_X1 _26771_ (.A(_08940_),
    .B1(_08799_),
    .B2(_08941_),
    .ZN(_02075_));
 AOI221_X2 _26772_ (.A(_03607_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .C1(_08869_),
    .C2(_10873_),
    .ZN(_08942_));
 NAND3_X1 _26773_ (.A1(_12935_),
    .A2(_13024_),
    .A3(_08929_),
    .ZN(_08943_));
 XNOR2_X1 _26774_ (.A(_00059_),
    .B(_08943_),
    .ZN(_08944_));
 AOI21_X2 _26775_ (.A(_08942_),
    .B1(_08944_),
    .B2(_08801_),
    .ZN(_08945_));
 AOI221_X2 _26776_ (.A(_08798_),
    .B1(_08939_),
    .B2(_08945_),
    .C1(_08595_),
    .C2(_07689_),
    .ZN(_08946_));
 INV_X1 _26777_ (.A(\cs_registers_i.mtval_q[25] ),
    .ZN(_08947_));
 AOI21_X1 _26778_ (.A(_08946_),
    .B1(_08799_),
    .B2(_08947_),
    .ZN(_02076_));
 NAND2_X2 _26779_ (.A1(_06989_),
    .A2(_08620_),
    .ZN(_08948_));
 NAND4_X1 _26780_ (.A1(_12935_),
    .A2(_13024_),
    .A3(\cs_registers_i.pc_id_i[25] ),
    .A4(_08935_),
    .ZN(_08949_));
 XNOR2_X1 _26781_ (.A(_00060_),
    .B(_08949_),
    .ZN(_08950_));
 AOI22_X1 _26782_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(_08792_),
    .B1(_08870_),
    .B2(_10874_),
    .ZN(_08951_));
 MUX2_X1 _26783_ (.A(_08950_),
    .B(_08951_),
    .S(_08854_),
    .Z(_08952_));
 OAI22_X2 _26784_ (.A1(_08163_),
    .A2(_08633_),
    .B1(_08948_),
    .B2(_08952_),
    .ZN(_08953_));
 MUX2_X1 _26785_ (.A(_08953_),
    .B(\cs_registers_i.mtval_q[26] ),
    .S(_08926_),
    .Z(_02077_));
 AND4_X1 _26786_ (.A1(_12935_),
    .A2(_13024_),
    .A3(\cs_registers_i.pc_id_i[25] ),
    .A4(\cs_registers_i.pc_id_i[26] ),
    .ZN(_08954_));
 NAND2_X1 _26787_ (.A1(_08929_),
    .A2(_08954_),
    .ZN(_08955_));
 XNOR2_X1 _26788_ (.A(_00061_),
    .B(_08955_),
    .ZN(_08956_));
 AOI22_X1 _26789_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(_08792_),
    .B1(_08870_),
    .B2(_10500_),
    .ZN(_08957_));
 MUX2_X1 _26790_ (.A(_08956_),
    .B(_08957_),
    .S(_08854_),
    .Z(_08958_));
 OAI22_X2 _26791_ (.A1(_07709_),
    .A2(_08633_),
    .B1(_08948_),
    .B2(_08958_),
    .ZN(_08959_));
 MUX2_X1 _26792_ (.A(_08959_),
    .B(\cs_registers_i.mtval_q[27] ),
    .S(_08926_),
    .Z(_02078_));
 AOI221_X2 _26793_ (.A(_03607_),
    .B1(_08791_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .C1(_08869_),
    .C2(net305),
    .ZN(_08960_));
 AND2_X1 _26794_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_08954_),
    .ZN(_08961_));
 NAND2_X1 _26795_ (.A1(_08935_),
    .A2(_08961_),
    .ZN(_08962_));
 XNOR2_X1 _26796_ (.A(_00062_),
    .B(_08962_),
    .ZN(_08963_));
 AOI21_X2 _26797_ (.A(_08960_),
    .B1(_08963_),
    .B2(_08801_),
    .ZN(_08964_));
 AOI221_X2 _26798_ (.A(_08798_),
    .B1(_08939_),
    .B2(_08964_),
    .C1(_08595_),
    .C2(_07718_),
    .ZN(_08965_));
 INV_X1 _26799_ (.A(\cs_registers_i.mtval_q[28] ),
    .ZN(_08966_));
 AOI21_X1 _26800_ (.A(_08965_),
    .B1(_08799_),
    .B2(_08966_),
    .ZN(_02079_));
 NAND3_X1 _26801_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_08929_),
    .A3(_08961_),
    .ZN(_08967_));
 XNOR2_X1 _26802_ (.A(_00063_),
    .B(_08967_),
    .ZN(_08968_));
 AOI22_X1 _26803_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(_08792_),
    .B1(_08870_),
    .B2(_10502_),
    .ZN(_08969_));
 MUX2_X1 _26804_ (.A(_08968_),
    .B(_08969_),
    .S(_08854_),
    .Z(_08970_));
 OAI22_X2 _26805_ (.A1(_07728_),
    .A2(_08633_),
    .B1(_08948_),
    .B2(_08970_),
    .ZN(_08971_));
 MUX2_X1 _26806_ (.A(_08971_),
    .B(\cs_registers_i.mtval_q[29] ),
    .S(_08926_),
    .Z(_02080_));
 MUX2_X2 _26807_ (.A(_00015_),
    .B(_00016_),
    .S(_08813_),
    .Z(_08972_));
 OAI221_X1 _26808_ (.A(_08599_),
    .B1(_08603_),
    .B2(_11435_),
    .C1(_08972_),
    .C2(_08815_),
    .ZN(_08973_));
 NOR2_X1 _26809_ (.A1(_00012_),
    .A2(_08803_),
    .ZN(_08974_));
 AOI21_X1 _26810_ (.A(_08974_),
    .B1(_15537_),
    .B2(_08803_),
    .ZN(_08975_));
 NAND2_X1 _26811_ (.A1(_08875_),
    .A2(_08975_),
    .ZN(_08976_));
 NAND4_X1 _26812_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08973_),
    .A4(_08976_),
    .ZN(_08977_));
 OAI21_X1 _26813_ (.A(_08977_),
    .B1(_08905_),
    .B2(_07492_),
    .ZN(_08978_));
 MUX2_X1 _26814_ (.A(_08978_),
    .B(\cs_registers_i.mtval_q[2] ),
    .S(_08926_),
    .Z(_02081_));
 AND3_X1 _26815_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(\cs_registers_i.pc_id_i[29] ),
    .A3(_08961_),
    .ZN(_08979_));
 NAND2_X1 _26816_ (.A1(_08935_),
    .A2(_08979_),
    .ZN(_08980_));
 XNOR2_X1 _26817_ (.A(_00064_),
    .B(_08980_),
    .ZN(_08981_));
 AOI22_X1 _26818_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(_08792_),
    .B1(_08870_),
    .B2(_10498_),
    .ZN(_08982_));
 MUX2_X1 _26819_ (.A(_08981_),
    .B(_08982_),
    .S(_08854_),
    .Z(_08983_));
 OAI22_X1 _26820_ (.A1(_07983_),
    .A2(_08633_),
    .B1(_08948_),
    .B2(_08983_),
    .ZN(_08984_));
 MUX2_X1 _26821_ (.A(_08984_),
    .B(\cs_registers_i.mtval_q[30] ),
    .S(_08926_),
    .Z(_02082_));
 AOI22_X1 _26822_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(_08792_),
    .B1(_08870_),
    .B2(_10509_),
    .ZN(_08985_));
 NAND2_X1 _26823_ (.A1(_08599_),
    .A2(_08985_),
    .ZN(_08986_));
 NAND3_X1 _26824_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(_08929_),
    .A3(_08979_),
    .ZN(_08987_));
 XOR2_X1 _26825_ (.A(_00065_),
    .B(_08987_),
    .Z(_08988_));
 OAI21_X1 _26826_ (.A(_08986_),
    .B1(_08988_),
    .B2(_08599_),
    .ZN(_08989_));
 OAI22_X1 _26827_ (.A1(_07748_),
    .A2(_08633_),
    .B1(_08948_),
    .B2(_08989_),
    .ZN(_08990_));
 MUX2_X1 _26828_ (.A(_08990_),
    .B(\cs_registers_i.mtval_q[31] ),
    .S(_08926_),
    .Z(_02083_));
 XNOR2_X1 _26829_ (.A(_00019_),
    .B(_08820_),
    .ZN(_08991_));
 NAND2_X1 _26830_ (.A1(_08802_),
    .A2(_08991_),
    .ZN(_08992_));
 INV_X1 _26831_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .ZN(_08993_));
 MUX2_X2 _26832_ (.A(_00017_),
    .B(_00018_),
    .S(_08813_),
    .Z(_08994_));
 OAI221_X1 _26833_ (.A(_08854_),
    .B1(_08603_),
    .B2(_08993_),
    .C1(_08994_),
    .C2(_08815_),
    .ZN(_08995_));
 NAND4_X1 _26834_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_08992_),
    .A4(_08995_),
    .ZN(_08996_));
 OAI21_X1 _26835_ (.A(_08996_),
    .B1(_08905_),
    .B2(_07791_),
    .ZN(_08997_));
 MUX2_X1 _26836_ (.A(_08997_),
    .B(\cs_registers_i.mtval_q[3] ),
    .S(_08926_),
    .Z(_02084_));
 NAND4_X1 _26837_ (.A1(_10675_),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(_11517_),
    .A4(_08803_),
    .ZN(_08998_));
 XNOR2_X1 _26838_ (.A(_00022_),
    .B(_08998_),
    .ZN(_08999_));
 NAND2_X1 _26839_ (.A1(_08802_),
    .A2(_08999_),
    .ZN(_09000_));
 MUX2_X2 _26840_ (.A(_00020_),
    .B(_00021_),
    .S(_08813_),
    .Z(_09001_));
 OAI221_X1 _26841_ (.A(_08854_),
    .B1(_08602_),
    .B2(_11556_),
    .C1(_09001_),
    .C2(_08815_),
    .ZN(_09002_));
 NAND4_X1 _26842_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_09000_),
    .A4(_09002_),
    .ZN(_09003_));
 OAI21_X1 _26843_ (.A(_09003_),
    .B1(_08905_),
    .B2(_07800_),
    .ZN(_09004_));
 MUX2_X1 _26844_ (.A(_09004_),
    .B(\cs_registers_i.mtval_q[4] ),
    .S(_08926_),
    .Z(_02085_));
 INV_X1 _26845_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .ZN(_09005_));
 MUX2_X2 _26846_ (.A(_00023_),
    .B(_00024_),
    .S(_10338_),
    .Z(_09006_));
 OAI221_X1 _26847_ (.A(_08598_),
    .B1(_08602_),
    .B2(_09005_),
    .C1(_09006_),
    .C2(_08601_),
    .ZN(_09007_));
 NAND4_X1 _26848_ (.A1(_11517_),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(_08803_),
    .A4(_15536_),
    .ZN(_09008_));
 XOR2_X1 _26849_ (.A(_00025_),
    .B(_09008_),
    .Z(_09009_));
 OAI21_X1 _26850_ (.A(_09007_),
    .B1(_09009_),
    .B2(_08598_),
    .ZN(_09010_));
 NOR2_X1 _26851_ (.A1(_08621_),
    .A2(_09010_),
    .ZN(_09011_));
 MUX2_X1 _26852_ (.A(_07810_),
    .B(_09011_),
    .S(_08620_),
    .Z(_09012_));
 MUX2_X1 _26853_ (.A(_09012_),
    .B(\cs_registers_i.mtval_q[5] ),
    .S(_08798_),
    .Z(_02086_));
 NOR2_X1 _26854_ (.A1(_08804_),
    .A2(_08805_),
    .ZN(_09013_));
 XOR2_X1 _26855_ (.A(_00027_),
    .B(_09013_),
    .Z(_09014_));
 NAND2_X1 _26856_ (.A1(_08802_),
    .A2(_09014_),
    .ZN(_09015_));
 INV_X1 _26857_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .ZN(_09016_));
 MUX2_X2 _26858_ (.A(_10301_),
    .B(_00026_),
    .S(_10338_),
    .Z(_09017_));
 OAI221_X1 _26859_ (.A(_08854_),
    .B1(_08602_),
    .B2(_09016_),
    .C1(_09017_),
    .C2(_08815_),
    .ZN(_09018_));
 NAND4_X1 _26860_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_09015_),
    .A4(_09018_),
    .ZN(_09019_));
 OAI21_X1 _26861_ (.A(_09019_),
    .B1(_08905_),
    .B2(_07821_),
    .ZN(_09020_));
 MUX2_X1 _26862_ (.A(_09020_),
    .B(\cs_registers_i.mtval_q[6] ),
    .S(_08798_),
    .Z(_02087_));
 NAND3_X1 _26863_ (.A1(_08803_),
    .A2(_15536_),
    .A3(_08806_),
    .ZN(_09021_));
 XNOR2_X1 _26864_ (.A(_00029_),
    .B(_09021_),
    .ZN(_09022_));
 NAND2_X1 _26865_ (.A1(_08802_),
    .A2(_09022_),
    .ZN(_09023_));
 INV_X1 _26866_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .ZN(_09024_));
 MUX2_X1 _26867_ (.A(_00216_),
    .B(_00028_),
    .S(_10338_),
    .Z(_09025_));
 OAI221_X1 _26868_ (.A(_08854_),
    .B1(_08602_),
    .B2(_09024_),
    .C1(_09025_),
    .C2(_08601_),
    .ZN(_09026_));
 NAND4_X1 _26869_ (.A1(_08597_),
    .A2(_08819_),
    .A3(_09023_),
    .A4(_09026_),
    .ZN(_09027_));
 OAI21_X1 _26870_ (.A(_09027_),
    .B1(_08905_),
    .B2(_07828_),
    .ZN(_09028_));
 MUX2_X1 _26871_ (.A(_09028_),
    .B(\cs_registers_i.mtval_q[7] ),
    .S(_08798_),
    .Z(_02088_));
 NAND2_X1 _26872_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(_08799_),
    .ZN(_09029_));
 INV_X1 _26873_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .ZN(_09030_));
 MUX2_X2 _26874_ (.A(_00030_),
    .B(_00031_),
    .S(_10338_),
    .Z(_09031_));
 OAI221_X2 _26875_ (.A(_08598_),
    .B1(_08602_),
    .B2(_09030_),
    .C1(_09031_),
    .C2(_08601_),
    .ZN(_09032_));
 XNOR2_X1 _26876_ (.A(_00032_),
    .B(_08808_),
    .ZN(_09033_));
 OAI21_X1 _26877_ (.A(_09032_),
    .B1(_09033_),
    .B2(_08599_),
    .ZN(_09034_));
 NOR3_X1 _26878_ (.A1(_08621_),
    .A2(_08596_),
    .A3(_09034_),
    .ZN(_09035_));
 AOI21_X1 _26879_ (.A(_09035_),
    .B1(_08757_),
    .B2(_07844_),
    .ZN(_09036_));
 OAI21_X1 _26880_ (.A(_09029_),
    .B1(_09036_),
    .B2(_08799_),
    .ZN(_02089_));
 INV_X1 _26881_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .ZN(_09037_));
 MUX2_X2 _26882_ (.A(_00033_),
    .B(_00034_),
    .S(_10338_),
    .Z(_09038_));
 OAI221_X1 _26883_ (.A(_08598_),
    .B1(_08602_),
    .B2(_09037_),
    .C1(_09038_),
    .C2(_08601_),
    .ZN(_09039_));
 NAND2_X1 _26884_ (.A1(_11788_),
    .A2(_08821_),
    .ZN(_09040_));
 XOR2_X2 _26885_ (.A(_00035_),
    .B(_09040_),
    .Z(_09041_));
 OAI21_X1 _26886_ (.A(_09039_),
    .B1(_09041_),
    .B2(_08598_),
    .ZN(_09042_));
 NOR2_X1 _26887_ (.A1(_08621_),
    .A2(_09042_),
    .ZN(_09043_));
 MUX2_X1 _26888_ (.A(_07854_),
    .B(_09043_),
    .S(_08620_),
    .Z(_09044_));
 MUX2_X1 _26889_ (.A(_09044_),
    .B(\cs_registers_i.mtval_q[9] ),
    .S(_08798_),
    .Z(_02090_));
 NAND2_X2 _26890_ (.A1(_05199_),
    .A2(_07488_),
    .ZN(_09045_));
 CLKBUF_X3 _26891_ (.A(_09045_),
    .Z(_09046_));
 NAND2_X1 _26892_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(_09046_),
    .ZN(_09047_));
 OAI21_X1 _26893_ (.A(_09047_),
    .B1(_09046_),
    .B2(_07525_),
    .ZN(_09048_));
 BUF_X4 _26894_ (.A(_03876_),
    .Z(_09049_));
 MUX2_X1 _26895_ (.A(net3),
    .B(_09048_),
    .S(_09049_),
    .Z(_02091_));
 CLKBUF_X3 _26896_ (.A(_09045_),
    .Z(_09050_));
 MUX2_X1 _26897_ (.A(_08275_),
    .B(\cs_registers_i.csr_mtvec_o[11] ),
    .S(_09050_),
    .Z(_09051_));
 MUX2_X1 _26898_ (.A(net4),
    .B(_09051_),
    .S(_09049_),
    .Z(_02092_));
 MUX2_X1 _26899_ (.A(_08444_),
    .B(\cs_registers_i.csr_mtvec_o[12] ),
    .S(_09050_),
    .Z(_09052_));
 MUX2_X1 _26900_ (.A(net5),
    .B(_09052_),
    .S(_09049_),
    .Z(_02093_));
 BUF_X4 _26901_ (.A(_09045_),
    .Z(_09053_));
 MUX2_X1 _26902_ (.A(_07569_),
    .B(\cs_registers_i.csr_mtvec_o[13] ),
    .S(_09053_),
    .Z(_09054_));
 MUX2_X1 _26903_ (.A(net6),
    .B(_09054_),
    .S(_09049_),
    .Z(_02094_));
 MUX2_X1 _26904_ (.A(_07579_),
    .B(\cs_registers_i.csr_mtvec_o[14] ),
    .S(_09053_),
    .Z(_09055_));
 MUX2_X1 _26905_ (.A(net7),
    .B(_09055_),
    .S(_09049_),
    .Z(_02095_));
 MUX2_X1 _26906_ (.A(_08299_),
    .B(\cs_registers_i.csr_mtvec_o[15] ),
    .S(_09053_),
    .Z(_09056_));
 MUX2_X1 _26907_ (.A(net8),
    .B(_09056_),
    .S(_09049_),
    .Z(_02096_));
 MUX2_X1 _26908_ (.A(_07600_),
    .B(\cs_registers_i.csr_mtvec_o[16] ),
    .S(_09053_),
    .Z(_09057_));
 MUX2_X1 _26909_ (.A(net9),
    .B(_09057_),
    .S(_09049_),
    .Z(_02097_));
 NAND2_X1 _26910_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(_09050_),
    .ZN(_09058_));
 OAI21_X1 _26911_ (.A(_09058_),
    .B1(_09046_),
    .B2(_08312_),
    .ZN(_09059_));
 MUX2_X1 _26912_ (.A(net10),
    .B(_09059_),
    .S(_09049_),
    .Z(_02098_));
 MUX2_X1 _26913_ (.A(_07914_),
    .B(\cs_registers_i.csr_mtvec_o[18] ),
    .S(_09053_),
    .Z(_09060_));
 MUX2_X1 _26914_ (.A(net11),
    .B(_09060_),
    .S(_09049_),
    .Z(_02099_));
 NAND2_X1 _26915_ (.A1(\cs_registers_i.csr_mtvec_o[19] ),
    .A2(_09050_),
    .ZN(_09061_));
 OAI21_X1 _26916_ (.A(_09061_),
    .B1(_09046_),
    .B2(_07624_),
    .ZN(_09062_));
 MUX2_X1 _26917_ (.A(net12),
    .B(_09062_),
    .S(_09049_),
    .Z(_02100_));
 NAND2_X1 _26918_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_09050_),
    .ZN(_09063_));
 OAI21_X1 _26919_ (.A(_09063_),
    .B1(_09046_),
    .B2(_07640_),
    .ZN(_09064_));
 CLKBUF_X3 _26920_ (.A(_03876_),
    .Z(_09065_));
 MUX2_X1 _26921_ (.A(net13),
    .B(_09064_),
    .S(_09065_),
    .Z(_02101_));
 MUX2_X1 _26922_ (.A(_08343_),
    .B(\cs_registers_i.csr_mtvec_o[21] ),
    .S(_09053_),
    .Z(_09066_));
 MUX2_X1 _26923_ (.A(net23),
    .B(_09066_),
    .S(_09065_),
    .Z(_02102_));
 NAND2_X1 _26924_ (.A1(\cs_registers_i.csr_mtvec_o[22] ),
    .A2(_09050_),
    .ZN(_09067_));
 OAI21_X1 _26925_ (.A(_09067_),
    .B1(_09046_),
    .B2(_07657_),
    .ZN(_09068_));
 MUX2_X1 _26926_ (.A(net24),
    .B(_09068_),
    .S(_09065_),
    .Z(_02103_));
 MUX2_X1 _26927_ (.A(_08355_),
    .B(\cs_registers_i.csr_mtvec_o[23] ),
    .S(_09053_),
    .Z(_09069_));
 MUX2_X1 _26928_ (.A(net25),
    .B(_09069_),
    .S(_09065_),
    .Z(_02104_));
 MUX2_X1 _26929_ (.A(_08149_),
    .B(\cs_registers_i.csr_mtvec_o[24] ),
    .S(_09053_),
    .Z(_09070_));
 MUX2_X1 _26930_ (.A(net26),
    .B(_09070_),
    .S(_09065_),
    .Z(_02105_));
 MUX2_X1 _26931_ (.A(_07689_),
    .B(\cs_registers_i.csr_mtvec_o[25] ),
    .S(_09053_),
    .Z(_09071_));
 MUX2_X1 _26932_ (.A(net27),
    .B(_09071_),
    .S(_09065_),
    .Z(_02106_));
 NAND2_X1 _26933_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(_09050_),
    .ZN(_09072_));
 OAI21_X1 _26934_ (.A(_09072_),
    .B1(_09046_),
    .B2(_08163_),
    .ZN(_09073_));
 MUX2_X1 _26935_ (.A(net28),
    .B(_09073_),
    .S(_09065_),
    .Z(_02107_));
 NAND2_X1 _26936_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_09050_),
    .ZN(_09074_));
 OAI21_X1 _26937_ (.A(_09074_),
    .B1(_09046_),
    .B2(_07709_),
    .ZN(_09075_));
 MUX2_X1 _26938_ (.A(net29),
    .B(_09075_),
    .S(_09065_),
    .Z(_02108_));
 MUX2_X1 _26939_ (.A(_07718_),
    .B(\cs_registers_i.csr_mtvec_o[28] ),
    .S(_09053_),
    .Z(_09076_));
 MUX2_X1 _26940_ (.A(net30),
    .B(_09076_),
    .S(_09065_),
    .Z(_02109_));
 NAND2_X1 _26941_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(_09050_),
    .ZN(_09077_));
 OAI21_X1 _26942_ (.A(_09077_),
    .B1(_09046_),
    .B2(_07728_),
    .ZN(_09078_));
 MUX2_X1 _26943_ (.A(net31),
    .B(_09078_),
    .S(_09065_),
    .Z(_02110_));
 NAND2_X1 _26944_ (.A1(\cs_registers_i.csr_mtvec_o[30] ),
    .A2(_09050_),
    .ZN(_09079_));
 OAI21_X1 _26945_ (.A(_09079_),
    .B1(_09046_),
    .B2(_07983_),
    .ZN(_09080_));
 MUX2_X1 _26946_ (.A(net32),
    .B(_09080_),
    .S(_03876_),
    .Z(_02111_));
 MUX2_X1 _26947_ (.A(_08405_),
    .B(\cs_registers_i.csr_mtvec_o[31] ),
    .S(_09045_),
    .Z(_09081_));
 MUX2_X1 _26948_ (.A(net33),
    .B(_09081_),
    .S(_03876_),
    .Z(_02112_));
 MUX2_X1 _26949_ (.A(_07844_),
    .B(\cs_registers_i.csr_mtvec_o[8] ),
    .S(_09045_),
    .Z(_09082_));
 MUX2_X1 _26950_ (.A(net34),
    .B(_09082_),
    .S(_03876_),
    .Z(_02113_));
 MUX2_X1 _26951_ (.A(_07854_),
    .B(\cs_registers_i.csr_mtvec_o[9] ),
    .S(_09045_),
    .Z(_09083_));
 MUX2_X1 _26952_ (.A(net35),
    .B(_09083_),
    .S(_03876_),
    .Z(_02114_));
 NAND3_X1 _26953_ (.A1(_03647_),
    .A2(_03451_),
    .A3(_06387_),
    .ZN(_09084_));
 MUX2_X1 _26954_ (.A(_03646_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .S(_09084_),
    .Z(_02115_));
 NAND2_X1 _26955_ (.A1(_06412_),
    .A2(_03615_),
    .ZN(_09085_));
 NOR4_X1 _26956_ (.A1(_03617_),
    .A2(_03647_),
    .A3(_03611_),
    .A4(_15538_),
    .ZN(_09086_));
 OAI21_X1 _26957_ (.A(_09085_),
    .B1(_09086_),
    .B2(_03615_),
    .ZN(_02116_));
 NOR3_X1 _26958_ (.A1(_03617_),
    .A2(_03647_),
    .A3(_03611_),
    .ZN(_09087_));
 NAND2_X1 _26959_ (.A1(_06421_),
    .A2(_09087_),
    .ZN(_09088_));
 MUX2_X1 _26960_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(_09088_),
    .S(_03451_),
    .Z(_02117_));
 NAND2_X1 _26961_ (.A1(_03445_),
    .A2(_03615_),
    .ZN(_09089_));
 NOR4_X1 _26962_ (.A1(_03617_),
    .A2(_03647_),
    .A3(_03611_),
    .A4(_06428_),
    .ZN(_09090_));
 OAI21_X1 _26963_ (.A(_09089_),
    .B1(_09090_),
    .B2(_03615_),
    .ZN(_02118_));
 NAND2_X1 _26964_ (.A1(_03444_),
    .A2(_03615_),
    .ZN(_09091_));
 NOR4_X1 _26965_ (.A1(_03617_),
    .A2(_03647_),
    .A3(_03611_),
    .A4(_06418_),
    .ZN(_09092_));
 OAI21_X1 _26966_ (.A(_09091_),
    .B1(_09092_),
    .B2(_03615_),
    .ZN(_02119_));
 NAND2_X1 _26967_ (.A1(_06446_),
    .A2(_09087_),
    .ZN(_09093_));
 MUX2_X1 _26968_ (.A(_06613_),
    .B(_09093_),
    .S(_03451_),
    .Z(_02120_));
 MUX2_X1 _26969_ (.A(_04045_),
    .B(\alu_adder_result_ex[0] ),
    .S(_03791_),
    .Z(_09094_));
 NOR2_X4 _26970_ (.A1(_04038_),
    .A2(_03441_),
    .ZN(_09095_));
 CLKBUF_X3 _26971_ (.A(_09095_),
    .Z(_09096_));
 MUX2_X1 _26972_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .B(_09094_),
    .S(_09096_),
    .Z(_02121_));
 MUX2_X1 _26973_ (.A(_11898_),
    .B(net386),
    .S(_03791_),
    .Z(_09097_));
 MUX2_X1 _26974_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .B(_09097_),
    .S(_09096_),
    .Z(_02122_));
 MUX2_X1 _26975_ (.A(_11398_),
    .B(\alu_adder_result_ex[11] ),
    .S(_03791_),
    .Z(_09098_));
 MUX2_X1 _26976_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .B(_09098_),
    .S(_09096_),
    .Z(_02123_));
 MUX2_X1 _26977_ (.A(_10868_),
    .B(\alu_adder_result_ex[12] ),
    .S(_03791_),
    .Z(_09099_));
 MUX2_X1 _26978_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .B(_09099_),
    .S(_09096_),
    .Z(_02124_));
 MUX2_X1 _26979_ (.A(_12075_),
    .B(\alu_adder_result_ex[13] ),
    .S(_03791_),
    .Z(_09100_));
 MUX2_X1 _26980_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .B(_09100_),
    .S(_09096_),
    .Z(_02125_));
 MUX2_X1 _26981_ (.A(_12177_),
    .B(net380),
    .S(_03791_),
    .Z(_09101_));
 MUX2_X1 _26982_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .B(_09101_),
    .S(_09096_),
    .Z(_02126_));
 MUX2_X1 _26983_ (.A(_12254_),
    .B(\alu_adder_result_ex[15] ),
    .S(_03791_),
    .Z(_09102_));
 MUX2_X1 _26984_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .B(_09102_),
    .S(_09096_),
    .Z(_02127_));
 MUX2_X1 _26985_ (.A(_12350_),
    .B(\alu_adder_result_ex[16] ),
    .S(_03791_),
    .Z(_09103_));
 MUX2_X1 _26986_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .B(_09103_),
    .S(_09096_),
    .Z(_02128_));
 MUX2_X1 _26987_ (.A(_12425_),
    .B(\alu_adder_result_ex[17] ),
    .S(_03791_),
    .Z(_09104_));
 CLKBUF_X3 _26988_ (.A(_09095_),
    .Z(_09105_));
 MUX2_X1 _26989_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .B(_09104_),
    .S(_09105_),
    .Z(_02129_));
 CLKBUF_X3 _26990_ (.A(_03790_),
    .Z(_09106_));
 MUX2_X1 _26991_ (.A(_12514_),
    .B(net371),
    .S(_09106_),
    .Z(_09107_));
 MUX2_X1 _26992_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .B(_09107_),
    .S(_09105_),
    .Z(_02130_));
 MUX2_X1 _26993_ (.A(_12589_),
    .B(net381),
    .S(_09106_),
    .Z(_09108_));
 MUX2_X1 _26994_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .B(_09108_),
    .S(_09105_),
    .Z(_02131_));
 MUX2_X1 _26995_ (.A(_03681_),
    .B(\alu_adder_result_ex[1] ),
    .S(_09106_),
    .Z(_09109_));
 MUX2_X1 _26996_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .B(_09109_),
    .S(_09105_),
    .Z(_02132_));
 MUX2_X1 _26997_ (.A(net359),
    .B(\alu_adder_result_ex[20] ),
    .S(_09106_),
    .Z(_09110_));
 MUX2_X1 _26998_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .B(_09110_),
    .S(_09105_),
    .Z(_02133_));
 MUX2_X1 _26999_ (.A(net361),
    .B(net366),
    .S(_09106_),
    .Z(_09111_));
 MUX2_X1 _27000_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .B(_09111_),
    .S(_09105_),
    .Z(_02134_));
 MUX2_X1 _27001_ (.A(_03713_),
    .B(\alu_adder_result_ex[22] ),
    .S(_09106_),
    .Z(_09112_));
 MUX2_X1 _27002_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .B(_09112_),
    .S(_09105_),
    .Z(_02135_));
 MUX2_X1 _27003_ (.A(_03724_),
    .B(net372),
    .S(_09106_),
    .Z(_09113_));
 MUX2_X1 _27004_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .B(_09113_),
    .S(_09105_),
    .Z(_02136_));
 MUX2_X1 _27005_ (.A(_03733_),
    .B(\alu_adder_result_ex[24] ),
    .S(_09106_),
    .Z(_09114_));
 MUX2_X1 _27006_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .B(_09114_),
    .S(_09105_),
    .Z(_02137_));
 MUX2_X1 _27007_ (.A(_13097_),
    .B(net373),
    .S(_09106_),
    .Z(_09115_));
 MUX2_X1 _27008_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .B(_09115_),
    .S(_09105_),
    .Z(_02138_));
 MUX2_X1 _27009_ (.A(net353),
    .B(net383),
    .S(_09106_),
    .Z(_09116_));
 CLKBUF_X3 _27010_ (.A(_09095_),
    .Z(_09117_));
 MUX2_X1 _27011_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .B(_09116_),
    .S(_09117_),
    .Z(_02139_));
 CLKBUF_X3 _27012_ (.A(_03790_),
    .Z(_09118_));
 MUX2_X1 _27013_ (.A(net343),
    .B(net376),
    .S(_09118_),
    .Z(_09119_));
 MUX2_X1 _27014_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B(_09119_),
    .S(_09117_),
    .Z(_02140_));
 MUX2_X1 _27015_ (.A(_03762_),
    .B(\alu_adder_result_ex[28] ),
    .S(_09118_),
    .Z(_09120_));
 MUX2_X1 _27016_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B(_09120_),
    .S(_09117_),
    .Z(_02141_));
 MUX2_X1 _27017_ (.A(_03769_),
    .B(net14),
    .S(_09118_),
    .Z(_09121_));
 MUX2_X1 _27018_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .B(_09121_),
    .S(_09117_),
    .Z(_02142_));
 MUX2_X1 _27019_ (.A(net295),
    .B(\alu_adder_result_ex[2] ),
    .S(_09118_),
    .Z(_09122_));
 MUX2_X1 _27020_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .B(_09122_),
    .S(_09117_),
    .Z(_02143_));
 MUX2_X1 _27021_ (.A(_03311_),
    .B(\alu_adder_result_ex[30] ),
    .S(_09118_),
    .Z(_09123_));
 MUX2_X1 _27022_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .B(_09123_),
    .S(_09117_),
    .Z(_02144_));
 OAI221_X1 _27023_ (.A(_09096_),
    .B1(_03789_),
    .B2(net279),
    .C1(_03371_),
    .C2(_03386_),
    .ZN(_09124_));
 OAI21_X1 _27024_ (.A(_09124_),
    .B1(_09096_),
    .B2(_06408_),
    .ZN(_02145_));
 MUX2_X1 _27025_ (.A(net320),
    .B(\alu_adder_result_ex[3] ),
    .S(_09118_),
    .Z(_09125_));
 MUX2_X1 _27026_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .B(_09125_),
    .S(_09117_),
    .Z(_02146_));
 MUX2_X1 _27027_ (.A(_11591_),
    .B(\alu_adder_result_ex[4] ),
    .S(_09118_),
    .Z(_09126_));
 MUX2_X1 _27028_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .B(_09126_),
    .S(_09117_),
    .Z(_02147_));
 MUX2_X1 _27029_ (.A(_11629_),
    .B(\alu_adder_result_ex[5] ),
    .S(_09118_),
    .Z(_09127_));
 MUX2_X1 _27030_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .B(_09127_),
    .S(_09117_),
    .Z(_02148_));
 MUX2_X1 _27031_ (.A(_11672_),
    .B(\alu_adder_result_ex[6] ),
    .S(_09118_),
    .Z(_09128_));
 MUX2_X1 _27032_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .B(_09128_),
    .S(_09117_),
    .Z(_02149_));
 MUX2_X1 _27033_ (.A(_03723_),
    .B(\alu_adder_result_ex[7] ),
    .S(_09118_),
    .Z(_09129_));
 MUX2_X1 _27034_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .B(_09129_),
    .S(_09095_),
    .Z(_02150_));
 MUX2_X1 _27035_ (.A(_03732_),
    .B(\alu_adder_result_ex[8] ),
    .S(_03790_),
    .Z(_09130_));
 MUX2_X1 _27036_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .B(_09130_),
    .S(_09095_),
    .Z(_02151_));
 MUX2_X1 _27037_ (.A(_11824_),
    .B(\alu_adder_result_ex[9] ),
    .S(_03790_),
    .Z(_09131_));
 MUX2_X1 _27038_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .B(_09131_),
    .S(_09095_),
    .Z(_02152_));
 OAI21_X2 _27039_ (.A(_03451_),
    .B1(_03617_),
    .B2(_03431_),
    .ZN(_09132_));
 CLKBUF_X3 _27040_ (.A(_09132_),
    .Z(_09133_));
 NAND2_X1 _27041_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .A2(_09133_),
    .ZN(_09134_));
 NAND2_X2 _27042_ (.A1(_03614_),
    .A2(_03451_),
    .ZN(_09135_));
 OAI21_X1 _27043_ (.A(_09134_),
    .B1(_09135_),
    .B2(_06402_),
    .ZN(_02153_));
 NOR2_X4 _27044_ (.A1(_03432_),
    .A2(_03441_),
    .ZN(_09136_));
 CLKBUF_X3 _27045_ (.A(_09136_),
    .Z(_09137_));
 AOI22_X1 _27046_ (.A1(_06551_),
    .A2(_09137_),
    .B1(_09133_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_09138_));
 INV_X1 _27047_ (.A(_09138_),
    .ZN(_02154_));
 NAND2_X1 _27048_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .A2(_09133_),
    .ZN(_09139_));
 INV_X1 _27049_ (.A(_00079_),
    .ZN(_09140_));
 INV_X1 _27050_ (.A(_06484_),
    .ZN(_09141_));
 AOI21_X1 _27051_ (.A(_09140_),
    .B1(_09141_),
    .B2(_06544_),
    .ZN(_09142_));
 OAI21_X1 _27052_ (.A(_09139_),
    .B1(_09135_),
    .B2(_09142_),
    .ZN(_02155_));
 AOI22_X1 _27053_ (.A1(_06571_),
    .A2(_09137_),
    .B1(_09133_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_09143_));
 INV_X1 _27054_ (.A(_09143_),
    .ZN(_02156_));
 AOI22_X1 _27055_ (.A1(_06581_),
    .A2(_09137_),
    .B1(_09133_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_09144_));
 INV_X1 _27056_ (.A(_09144_),
    .ZN(_02157_));
 CLKBUF_X3 _27057_ (.A(_09132_),
    .Z(_09145_));
 AOI22_X1 _27058_ (.A1(_06591_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_09146_));
 INV_X1 _27059_ (.A(_09146_),
    .ZN(_02158_));
 AOI22_X1 _27060_ (.A1(_06601_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .ZN(_09147_));
 INV_X1 _27061_ (.A(_09147_),
    .ZN(_02159_));
 NAND2_X1 _27062_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .A2(_09133_),
    .ZN(_09148_));
 OAI21_X1 _27063_ (.A(_09148_),
    .B1(_09135_),
    .B2(_06615_),
    .ZN(_02160_));
 AOI22_X1 _27064_ (.A1(_06622_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .ZN(_09149_));
 INV_X1 _27065_ (.A(_09149_),
    .ZN(_02161_));
 AOI22_X1 _27066_ (.A1(_06631_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .ZN(_09150_));
 INV_X1 _27067_ (.A(_09150_),
    .ZN(_02162_));
 AOI22_X1 _27068_ (.A1(_06640_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .ZN(_09151_));
 INV_X1 _27069_ (.A(_09151_),
    .ZN(_02163_));
 NAND2_X1 _27070_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .A2(_09133_),
    .ZN(_09152_));
 OAI21_X1 _27071_ (.A(_09152_),
    .B1(_09135_),
    .B2(_06462_),
    .ZN(_02164_));
 AOI22_X1 _27072_ (.A1(_06648_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .ZN(_09153_));
 INV_X1 _27073_ (.A(_09153_),
    .ZN(_02165_));
 AOI22_X1 _27074_ (.A1(_06658_),
    .A2(_09137_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .ZN(_09154_));
 INV_X1 _27075_ (.A(_09154_),
    .ZN(_02166_));
 CLKBUF_X3 _27076_ (.A(_09136_),
    .Z(_09155_));
 AOI22_X1 _27077_ (.A1(_06665_),
    .A2(_09155_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .ZN(_09156_));
 INV_X1 _27078_ (.A(_09156_),
    .ZN(_02167_));
 AOI22_X1 _27079_ (.A1(_06674_),
    .A2(_09155_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .ZN(_09157_));
 INV_X1 _27080_ (.A(_09157_),
    .ZN(_02168_));
 AOI22_X1 _27081_ (.A1(_06683_),
    .A2(_09155_),
    .B1(_09145_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .ZN(_09158_));
 INV_X1 _27082_ (.A(_09158_),
    .ZN(_02169_));
 CLKBUF_X3 _27083_ (.A(_09132_),
    .Z(_09159_));
 AOI22_X1 _27084_ (.A1(_06692_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .ZN(_09160_));
 INV_X1 _27085_ (.A(_09160_),
    .ZN(_02170_));
 AOI22_X1 _27086_ (.A1(_06702_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .ZN(_09161_));
 INV_X1 _27087_ (.A(_09161_),
    .ZN(_02171_));
 AOI21_X1 _27088_ (.A(_09135_),
    .B1(_06711_),
    .B2(_00095_),
    .ZN(_09162_));
 AOI21_X1 _27089_ (.A(_09162_),
    .B1(_09133_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .ZN(_09163_));
 INV_X1 _27090_ (.A(_09163_),
    .ZN(_02172_));
 NAND2_X1 _27091_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .A2(_09133_),
    .ZN(_09164_));
 OAI21_X1 _27092_ (.A(_09164_),
    .B1(_09135_),
    .B2(_06726_),
    .ZN(_02173_));
 AOI22_X1 _27093_ (.A1(_06733_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .ZN(_09165_));
 INV_X1 _27094_ (.A(_09165_),
    .ZN(_02174_));
 AOI22_X1 _27095_ (.A1(_06471_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_09166_));
 INV_X1 _27096_ (.A(_09166_),
    .ZN(_02175_));
 AOI22_X1 _27097_ (.A1(_06741_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_09167_));
 INV_X1 _27098_ (.A(_09167_),
    .ZN(_02176_));
 AOI22_X1 _27099_ (.A1(_06751_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .ZN(_09168_));
 INV_X1 _27100_ (.A(_09168_),
    .ZN(_02177_));
 AOI22_X1 _27101_ (.A1(_06485_),
    .A2(_09155_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_09169_));
 INV_X1 _27102_ (.A(_09169_),
    .ZN(_02178_));
 AOI22_X1 _27103_ (.A1(_06496_),
    .A2(_09136_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .ZN(_09170_));
 INV_X1 _27104_ (.A(_09170_),
    .ZN(_02179_));
 AOI22_X1 _27105_ (.A1(_06506_),
    .A2(_09136_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .ZN(_09171_));
 INV_X1 _27106_ (.A(_09171_),
    .ZN(_02180_));
 AOI22_X1 _27107_ (.A1(_06515_),
    .A2(_09136_),
    .B1(_09159_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .ZN(_09172_));
 INV_X1 _27108_ (.A(_09172_),
    .ZN(_02181_));
 AOI22_X1 _27109_ (.A1(_06523_),
    .A2(_09136_),
    .B1(_09132_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .ZN(_09173_));
 INV_X1 _27110_ (.A(_09173_),
    .ZN(_02182_));
 AOI22_X1 _27111_ (.A1(_06532_),
    .A2(_09136_),
    .B1(_09132_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_09174_));
 INV_X1 _27112_ (.A(_09174_),
    .ZN(_02183_));
 NAND2_X1 _27113_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .A2(_09133_),
    .ZN(_09175_));
 OAI21_X1 _27114_ (.A(_09175_),
    .B1(_09135_),
    .B2(_06545_),
    .ZN(_02184_));
 OR2_X1 _27115_ (.A1(fetch_enable_q),
    .A2(net70),
    .ZN(_02185_));
 AND2_X2 _27116_ (.A1(_05805_),
    .A2(_06245_),
    .ZN(_09176_));
 BUF_X4 _27117_ (.A(_09176_),
    .Z(_09177_));
 MUX2_X1 _27118_ (.A(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B(_06223_),
    .S(_09177_),
    .Z(_02186_));
 BUF_X2 _27119_ (.A(_05543_),
    .Z(_09178_));
 MUX2_X1 _27120_ (.A(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .B(_09178_),
    .S(_06229_),
    .Z(_02187_));
 BUF_X2 _27121_ (.A(_05579_),
    .Z(_09179_));
 MUX2_X1 _27122_ (.A(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .B(_09179_),
    .S(_06229_),
    .Z(_02188_));
 BUF_X2 _27123_ (.A(_05613_),
    .Z(_09180_));
 MUX2_X1 _27124_ (.A(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .B(_09180_),
    .S(_06229_),
    .Z(_02189_));
 BUF_X2 _27125_ (.A(_05652_),
    .Z(_09181_));
 MUX2_X1 _27126_ (.A(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .B(_09181_),
    .S(_06229_),
    .Z(_02190_));
 NAND2_X1 _27127_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .A2(_06240_),
    .ZN(_09182_));
 OAI21_X1 _27128_ (.A(_09182_),
    .B1(_06241_),
    .B2(_06222_),
    .ZN(_02191_));
 BUF_X2 _27129_ (.A(_05720_),
    .Z(_09183_));
 BUF_X4 _27130_ (.A(_06228_),
    .Z(_09184_));
 MUX2_X1 _27131_ (.A(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .B(_09183_),
    .S(_09184_),
    .Z(_02192_));
 BUF_X2 _27132_ (.A(_05761_),
    .Z(_09185_));
 MUX2_X1 _27133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .B(_09185_),
    .S(_09184_),
    .Z(_02193_));
 BUF_X2 _27134_ (.A(_05801_),
    .Z(_09186_));
 MUX2_X1 _27135_ (.A(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .B(_09186_),
    .S(_09184_),
    .Z(_02194_));
 NOR2_X1 _27136_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .A2(_06229_),
    .ZN(_09187_));
 AOI21_X1 _27137_ (.A(_09187_),
    .B1(_06229_),
    .B2(_05850_),
    .ZN(_02195_));
 BUF_X2 _27138_ (.A(_05889_),
    .Z(_09188_));
 MUX2_X1 _27139_ (.A(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .B(_09188_),
    .S(_09184_),
    .Z(_02196_));
 MUX2_X1 _27140_ (.A(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .B(_09185_),
    .S(_09177_),
    .Z(_02197_));
 BUF_X2 _27141_ (.A(_05927_),
    .Z(_09189_));
 MUX2_X1 _27142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .B(_09189_),
    .S(_09184_),
    .Z(_02198_));
 BUF_X4 _27143_ (.A(_05973_),
    .Z(_09190_));
 MUX2_X1 _27144_ (.A(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .B(_09190_),
    .S(_09184_),
    .Z(_02199_));
 NOR2_X1 _27145_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .A2(_06229_),
    .ZN(_09191_));
 AOI21_X1 _27146_ (.A(_09191_),
    .B1(_06229_),
    .B2(_06016_),
    .ZN(_02200_));
 BUF_X2 _27147_ (.A(_06061_),
    .Z(_09192_));
 MUX2_X1 _27148_ (.A(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .B(_09192_),
    .S(_09184_),
    .Z(_02201_));
 BUF_X2 _27149_ (.A(_06099_),
    .Z(_09193_));
 MUX2_X1 _27150_ (.A(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .B(_09193_),
    .S(_09184_),
    .Z(_02202_));
 NAND2_X1 _27151_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .A2(_06240_),
    .ZN(_09194_));
 OAI21_X1 _27152_ (.A(_09194_),
    .B1(_06241_),
    .B2(_06138_),
    .ZN(_02203_));
 BUF_X4 _27153_ (.A(_06173_),
    .Z(_09195_));
 MUX2_X1 _27154_ (.A(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .B(net404),
    .S(_09184_),
    .Z(_02204_));
 BUF_X2 _27155_ (.A(_06206_),
    .Z(_09196_));
 MUX2_X1 _27156_ (.A(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .B(_09196_),
    .S(_09184_),
    .Z(_02205_));
 BUF_X4 _27157_ (.A(_04601_),
    .Z(_09197_));
 MUX2_X1 _27158_ (.A(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .B(_09197_),
    .S(_06228_),
    .Z(_02206_));
 BUF_X2 _27159_ (.A(_04765_),
    .Z(_09198_));
 MUX2_X1 _27160_ (.A(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .B(_09198_),
    .S(_06228_),
    .Z(_02207_));
 MUX2_X1 _27161_ (.A(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B(_09186_),
    .S(_09177_),
    .Z(_02208_));
 NAND2_X1 _27162_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A2(_06240_),
    .ZN(_09199_));
 OAI21_X1 _27163_ (.A(_09199_),
    .B1(_06241_),
    .B2(_04908_),
    .ZN(_02209_));
 NAND2_X1 _27164_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A2(_06240_),
    .ZN(_09200_));
 OAI21_X4 _27165_ (.A(_09200_),
    .B1(_04978_),
    .B2(_06241_),
    .ZN(_02210_));
 BUF_X4 _27166_ (.A(_05036_),
    .Z(_09201_));
 MUX2_X1 _27167_ (.A(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .B(_09201_),
    .S(_06228_),
    .Z(_02211_));
 BUF_X4 _27168_ (.A(_04849_),
    .Z(_09202_));
 MUX2_X1 _27169_ (.A(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .B(net331),
    .S(_06228_),
    .Z(_02212_));
 MUX2_X1 _27170_ (.A(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .B(net408),
    .S(_06228_),
    .Z(_02213_));
 NAND2_X1 _27171_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A2(_06240_),
    .ZN(_09203_));
 OAI21_X4 _27172_ (.A(_09203_),
    .B1(_05148_),
    .B2(_06241_),
    .ZN(_02214_));
 MUX2_X1 _27173_ (.A(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .B(net392),
    .S(_06228_),
    .Z(_02215_));
 NAND2_X1 _27174_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A2(_06240_),
    .ZN(_09204_));
 OAI21_X4 _27175_ (.A(_09204_),
    .B1(net441),
    .B2(_06241_),
    .ZN(_02216_));
 AND3_X1 _27176_ (.A1(_05412_),
    .A2(_06225_),
    .A3(_06245_),
    .ZN(_09205_));
 BUF_X4 _27177_ (.A(_09205_),
    .Z(_09206_));
 BUF_X4 _27178_ (.A(_09206_),
    .Z(_09207_));
 MUX2_X1 _27179_ (.A(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .B(_06223_),
    .S(_09207_),
    .Z(_02217_));
 MUX2_X1 _27180_ (.A(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .B(_06236_),
    .S(_09207_),
    .Z(_02218_));
 NOR2_X1 _27181_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A2(_09177_),
    .ZN(_09208_));
 AOI21_X1 _27182_ (.A(_09208_),
    .B1(_09177_),
    .B2(_05850_),
    .ZN(_02219_));
 NAND3_X4 _27183_ (.A1(_06224_),
    .A2(_06226_),
    .A3(_06245_),
    .ZN(_09209_));
 BUF_X4 _27184_ (.A(_09209_),
    .Z(_09210_));
 NAND2_X1 _27185_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .A2(_09210_),
    .ZN(_09211_));
 OAI21_X1 _27186_ (.A(_09211_),
    .B1(_09210_),
    .B2(_05464_),
    .ZN(_02220_));
 NAND2_X1 _27187_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .A2(_09210_),
    .ZN(_09212_));
 OAI21_X1 _27188_ (.A(_09212_),
    .B1(_09210_),
    .B2(_05510_),
    .ZN(_02221_));
 MUX2_X1 _27189_ (.A(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .B(_09178_),
    .S(_09207_),
    .Z(_02222_));
 MUX2_X1 _27190_ (.A(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .B(_09179_),
    .S(_09207_),
    .Z(_02223_));
 BUF_X4 _27191_ (.A(_09206_),
    .Z(_09213_));
 MUX2_X1 _27192_ (.A(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .B(_09180_),
    .S(_09213_),
    .Z(_02224_));
 MUX2_X1 _27193_ (.A(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .B(_09181_),
    .S(_09213_),
    .Z(_02225_));
 NOR2_X1 _27194_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .A2(_09207_),
    .ZN(_09214_));
 AOI21_X1 _27195_ (.A(_09214_),
    .B1(_09207_),
    .B2(_05688_),
    .ZN(_02226_));
 MUX2_X1 _27196_ (.A(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .B(_09183_),
    .S(_09213_),
    .Z(_02227_));
 MUX2_X1 _27197_ (.A(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .B(_09185_),
    .S(_09213_),
    .Z(_02228_));
 MUX2_X1 _27198_ (.A(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .B(_09186_),
    .S(_09213_),
    .Z(_02229_));
 MUX2_X1 _27199_ (.A(_05890_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .S(_06246_),
    .Z(_02230_));
 NOR2_X1 _27200_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .A2(_09207_),
    .ZN(_09215_));
 AOI21_X1 _27201_ (.A(_09215_),
    .B1(_09207_),
    .B2(_05850_),
    .ZN(_02231_));
 MUX2_X1 _27202_ (.A(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .B(_09188_),
    .S(_09213_),
    .Z(_02232_));
 MUX2_X1 _27203_ (.A(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .B(_09189_),
    .S(_09213_),
    .Z(_02233_));
 MUX2_X1 _27204_ (.A(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .B(_09190_),
    .S(_09213_),
    .Z(_02234_));
 NOR2_X1 _27205_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .A2(_09207_),
    .ZN(_09216_));
 AOI21_X1 _27206_ (.A(_09216_),
    .B1(_09207_),
    .B2(_06016_),
    .ZN(_02235_));
 MUX2_X1 _27207_ (.A(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .B(_09192_),
    .S(_09213_),
    .Z(_02236_));
 MUX2_X1 _27208_ (.A(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .B(_09193_),
    .S(_09213_),
    .Z(_02237_));
 NAND2_X1 _27209_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .A2(_09210_),
    .ZN(_09217_));
 OAI21_X1 _27210_ (.A(_09217_),
    .B1(_09210_),
    .B2(_06138_),
    .ZN(_02238_));
 MUX2_X1 _27211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .B(net404),
    .S(_09206_),
    .Z(_02239_));
 MUX2_X1 _27212_ (.A(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .B(_09196_),
    .S(_09206_),
    .Z(_02240_));
 MUX2_X1 _27213_ (.A(_05928_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .S(_06246_),
    .Z(_02241_));
 MUX2_X1 _27214_ (.A(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .B(_09197_),
    .S(_09206_),
    .Z(_02242_));
 MUX2_X1 _27215_ (.A(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .B(_09198_),
    .S(_09206_),
    .Z(_02243_));
 NAND2_X1 _27216_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .A2(_09209_),
    .ZN(_09218_));
 OAI21_X1 _27217_ (.A(_09218_),
    .B1(_09210_),
    .B2(_04908_),
    .ZN(_02244_));
 NAND2_X1 _27218_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .A2(_09209_),
    .ZN(_09219_));
 OAI21_X4 _27219_ (.A(_09219_),
    .B1(_04978_),
    .B2(_09210_),
    .ZN(_02245_));
 MUX2_X1 _27220_ (.A(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .B(net419),
    .S(_09206_),
    .Z(_02246_));
 MUX2_X1 _27221_ (.A(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .B(_09202_),
    .S(_09206_),
    .Z(_02247_));
 MUX2_X1 _27222_ (.A(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .B(net408),
    .S(_09206_),
    .Z(_02248_));
 NAND2_X1 _27223_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .A2(_09209_),
    .ZN(_09220_));
 OAI21_X4 _27224_ (.A(_09220_),
    .B1(_05148_),
    .B2(_09210_),
    .ZN(_02249_));
 MUX2_X1 _27225_ (.A(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .B(net392),
    .S(_09206_),
    .Z(_02250_));
 NAND2_X1 _27226_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(_09209_),
    .ZN(_09221_));
 OAI21_X4 _27227_ (.A(_09221_),
    .B1(_05260_),
    .B2(_09210_),
    .ZN(_02251_));
 MUX2_X1 _27228_ (.A(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B(_09190_),
    .S(_09177_),
    .Z(_02252_));
 NOR2_X2 _27229_ (.A1(_10395_),
    .A2(_10902_),
    .ZN(_09222_));
 AND4_X1 _27230_ (.A1(_05412_),
    .A2(_04603_),
    .A3(_06225_),
    .A4(_09222_),
    .ZN(_09223_));
 BUF_X4 _27231_ (.A(_09223_),
    .Z(_09224_));
 BUF_X4 _27232_ (.A(_09224_),
    .Z(_09225_));
 MUX2_X1 _27233_ (.A(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .B(_06223_),
    .S(_09225_),
    .Z(_02253_));
 MUX2_X1 _27234_ (.A(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .B(_06236_),
    .S(_09225_),
    .Z(_02254_));
 NAND4_X4 _27235_ (.A1(_06224_),
    .A2(_04603_),
    .A3(_06226_),
    .A4(_09222_),
    .ZN(_09226_));
 CLKBUF_X3 _27236_ (.A(_09226_),
    .Z(_09227_));
 NAND2_X1 _27237_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .A2(_09227_),
    .ZN(_09228_));
 OAI21_X1 _27238_ (.A(_09228_),
    .B1(_09227_),
    .B2(_05464_),
    .ZN(_02255_));
 NAND2_X1 _27239_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .A2(_09227_),
    .ZN(_09229_));
 OAI21_X1 _27240_ (.A(_09229_),
    .B1(_09227_),
    .B2(_05510_),
    .ZN(_02256_));
 MUX2_X1 _27241_ (.A(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .B(_09178_),
    .S(_09225_),
    .Z(_02257_));
 MUX2_X1 _27242_ (.A(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .B(_09179_),
    .S(_09225_),
    .Z(_02258_));
 BUF_X4 _27243_ (.A(_09224_),
    .Z(_09230_));
 MUX2_X1 _27244_ (.A(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .B(_09180_),
    .S(_09230_),
    .Z(_02259_));
 MUX2_X1 _27245_ (.A(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .B(_09181_),
    .S(_09230_),
    .Z(_02260_));
 NOR2_X1 _27246_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .A2(_09225_),
    .ZN(_09231_));
 AOI21_X1 _27247_ (.A(_09231_),
    .B1(_09225_),
    .B2(_05688_),
    .ZN(_02261_));
 MUX2_X1 _27248_ (.A(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .B(_09183_),
    .S(_09230_),
    .Z(_02262_));
 NOR2_X1 _27249_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .A2(_09177_),
    .ZN(_09232_));
 AOI21_X1 _27250_ (.A(_09232_),
    .B1(_09177_),
    .B2(_06016_),
    .ZN(_02263_));
 MUX2_X1 _27251_ (.A(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .B(_09185_),
    .S(_09230_),
    .Z(_02264_));
 MUX2_X1 _27252_ (.A(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .B(_09186_),
    .S(_09230_),
    .Z(_02265_));
 NOR2_X1 _27253_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .A2(_09225_),
    .ZN(_09233_));
 AOI21_X1 _27254_ (.A(_09233_),
    .B1(_09225_),
    .B2(_05850_),
    .ZN(_02266_));
 MUX2_X1 _27255_ (.A(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .B(_09188_),
    .S(_09230_),
    .Z(_02267_));
 MUX2_X1 _27256_ (.A(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .B(_09189_),
    .S(_09230_),
    .Z(_02268_));
 MUX2_X1 _27257_ (.A(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .B(_09190_),
    .S(_09230_),
    .Z(_02269_));
 NOR2_X1 _27258_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .A2(_09225_),
    .ZN(_09234_));
 AOI21_X1 _27259_ (.A(_09234_),
    .B1(_09225_),
    .B2(_06016_),
    .ZN(_02270_));
 MUX2_X1 _27260_ (.A(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .B(_09192_),
    .S(_09230_),
    .Z(_02271_));
 MUX2_X1 _27261_ (.A(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .B(_09193_),
    .S(_09230_),
    .Z(_02272_));
 NAND2_X1 _27262_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .A2(_09227_),
    .ZN(_09235_));
 OAI21_X1 _27263_ (.A(_09235_),
    .B1(_09227_),
    .B2(_06138_),
    .ZN(_02273_));
 BUF_X4 _27264_ (.A(_09176_),
    .Z(_09236_));
 MUX2_X1 _27265_ (.A(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .B(_09192_),
    .S(_09236_),
    .Z(_02274_));
 MUX2_X1 _27266_ (.A(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .B(net404),
    .S(_09224_),
    .Z(_02275_));
 MUX2_X1 _27267_ (.A(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .B(_09196_),
    .S(_09224_),
    .Z(_02276_));
 MUX2_X1 _27268_ (.A(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .B(_09197_),
    .S(_09224_),
    .Z(_02277_));
 MUX2_X1 _27269_ (.A(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .B(_09198_),
    .S(_09224_),
    .Z(_02278_));
 NAND2_X1 _27270_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .A2(_09226_),
    .ZN(_09237_));
 OAI21_X1 _27271_ (.A(_09237_),
    .B1(_09227_),
    .B2(_04908_),
    .ZN(_02279_));
 NAND2_X1 _27272_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .A2(_09226_),
    .ZN(_09238_));
 OAI21_X4 _27273_ (.A(_09238_),
    .B1(net442),
    .B2(_09227_),
    .ZN(_02280_));
 MUX2_X1 _27274_ (.A(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .B(_09201_),
    .S(_09224_),
    .Z(_02281_));
 MUX2_X1 _27275_ (.A(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .B(_09202_),
    .S(_09224_),
    .Z(_02282_));
 MUX2_X1 _27276_ (.A(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .B(_05411_),
    .S(_09224_),
    .Z(_02283_));
 NAND2_X1 _27277_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A2(_09226_),
    .ZN(_09239_));
 OAI21_X4 _27278_ (.A(_09239_),
    .B1(net445),
    .B2(_09227_),
    .ZN(_02284_));
 MUX2_X1 _27279_ (.A(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B(_09193_),
    .S(_09236_),
    .Z(_02285_));
 MUX2_X1 _27280_ (.A(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .B(net392),
    .S(_09224_),
    .Z(_02286_));
 NAND2_X1 _27281_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A2(_09226_),
    .ZN(_09240_));
 OAI21_X4 _27282_ (.A(_09240_),
    .B1(_05260_),
    .B2(_09227_),
    .ZN(_02287_));
 AND3_X1 _27283_ (.A1(_05412_),
    .A2(_04852_),
    .A3(_06225_),
    .ZN(_09241_));
 BUF_X4 _27284_ (.A(_09241_),
    .Z(_09242_));
 BUF_X4 _27285_ (.A(_09242_),
    .Z(_09243_));
 MUX2_X1 _27286_ (.A(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .B(_06223_),
    .S(_09243_),
    .Z(_02288_));
 MUX2_X1 _27287_ (.A(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .B(_06236_),
    .S(_09243_),
    .Z(_02289_));
 NAND3_X4 _27288_ (.A1(_06224_),
    .A2(_04852_),
    .A3(_06226_),
    .ZN(_09244_));
 BUF_X4 _27289_ (.A(_09244_),
    .Z(_09245_));
 NAND2_X1 _27290_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .A2(_09245_),
    .ZN(_09246_));
 OAI21_X1 _27291_ (.A(_09246_),
    .B1(_09245_),
    .B2(_05464_),
    .ZN(_02290_));
 NAND2_X1 _27292_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .A2(_09245_),
    .ZN(_09247_));
 OAI21_X1 _27293_ (.A(_09247_),
    .B1(_09245_),
    .B2(_05510_),
    .ZN(_02291_));
 MUX2_X1 _27294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .B(_09178_),
    .S(_09243_),
    .Z(_02292_));
 MUX2_X1 _27295_ (.A(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .B(_09179_),
    .S(_09243_),
    .Z(_02293_));
 BUF_X4 _27296_ (.A(_09242_),
    .Z(_09248_));
 MUX2_X1 _27297_ (.A(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .B(_09180_),
    .S(_09248_),
    .Z(_02294_));
 MUX2_X1 _27298_ (.A(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .B(_09181_),
    .S(_09248_),
    .Z(_02295_));
 CLKBUF_X3 _27299_ (.A(_06246_),
    .Z(_09249_));
 NAND2_X1 _27300_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A2(_09249_),
    .ZN(_09250_));
 NAND2_X2 _27301_ (.A1(_05805_),
    .A2(_06245_),
    .ZN(_09251_));
 OAI21_X1 _27302_ (.A(_09250_),
    .B1(_09251_),
    .B2(_06138_),
    .ZN(_02296_));
 MUX2_X1 _27303_ (.A(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .B(_06236_),
    .S(_09236_),
    .Z(_02297_));
 NOR2_X1 _27304_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .A2(_09243_),
    .ZN(_09252_));
 AOI21_X1 _27305_ (.A(_09252_),
    .B1(_09243_),
    .B2(_05688_),
    .ZN(_02298_));
 MUX2_X1 _27306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .B(_09183_),
    .S(_09248_),
    .Z(_02299_));
 MUX2_X1 _27307_ (.A(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .B(_09185_),
    .S(_09248_),
    .Z(_02300_));
 MUX2_X1 _27308_ (.A(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .B(_09186_),
    .S(_09248_),
    .Z(_02301_));
 NOR2_X1 _27309_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .A2(_09243_),
    .ZN(_09253_));
 AOI21_X1 _27310_ (.A(_09253_),
    .B1(_09243_),
    .B2(_05850_),
    .ZN(_02302_));
 MUX2_X1 _27311_ (.A(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .B(_09188_),
    .S(_09248_),
    .Z(_02303_));
 MUX2_X1 _27312_ (.A(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .B(_09189_),
    .S(_09248_),
    .Z(_02304_));
 MUX2_X1 _27313_ (.A(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .B(_09190_),
    .S(_09248_),
    .Z(_02305_));
 NOR2_X1 _27314_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .A2(_09243_),
    .ZN(_09254_));
 AOI21_X1 _27315_ (.A(_09254_),
    .B1(_09243_),
    .B2(_06016_),
    .ZN(_02306_));
 MUX2_X1 _27316_ (.A(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .B(_09192_),
    .S(_09248_),
    .Z(_02307_));
 MUX2_X1 _27317_ (.A(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B(_09195_),
    .S(_09236_),
    .Z(_02308_));
 MUX2_X1 _27318_ (.A(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .B(_09193_),
    .S(_09248_),
    .Z(_02309_));
 NAND2_X1 _27319_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .A2(_09245_),
    .ZN(_09255_));
 OAI21_X1 _27320_ (.A(_09255_),
    .B1(_09245_),
    .B2(_06138_),
    .ZN(_02310_));
 MUX2_X1 _27321_ (.A(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .B(net404),
    .S(_09242_),
    .Z(_02311_));
 MUX2_X1 _27322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .B(_09196_),
    .S(_09242_),
    .Z(_02312_));
 MUX2_X1 _27323_ (.A(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .B(_09197_),
    .S(_09242_),
    .Z(_02313_));
 MUX2_X1 _27324_ (.A(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .B(_09198_),
    .S(_09242_),
    .Z(_02314_));
 NAND2_X1 _27325_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .A2(_09244_),
    .ZN(_09256_));
 OAI21_X1 _27326_ (.A(_09256_),
    .B1(_09245_),
    .B2(_04908_),
    .ZN(_02315_));
 NAND2_X1 _27327_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .A2(_09244_),
    .ZN(_09257_));
 OAI21_X1 _27328_ (.A(_09257_),
    .B1(_09245_),
    .B2(_04978_),
    .ZN(_02316_));
 MUX2_X1 _27329_ (.A(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .B(net419),
    .S(_09242_),
    .Z(_02317_));
 MUX2_X1 _27330_ (.A(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .B(net331),
    .S(_09242_),
    .Z(_02318_));
 MUX2_X1 _27331_ (.A(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .B(_09196_),
    .S(_09236_),
    .Z(_02319_));
 MUX2_X1 _27332_ (.A(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .B(net408),
    .S(_09242_),
    .Z(_02320_));
 NAND2_X1 _27333_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .A2(_09244_),
    .ZN(_09258_));
 OAI21_X4 _27334_ (.A(_09258_),
    .B1(_05148_),
    .B2(_09245_),
    .ZN(_02321_));
 MUX2_X1 _27335_ (.A(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .B(_06208_),
    .S(_09242_),
    .Z(_02322_));
 NAND2_X1 _27336_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .A2(_09244_),
    .ZN(_09259_));
 OAI21_X4 _27337_ (.A(_09259_),
    .B1(_05260_),
    .B2(_09245_),
    .ZN(_02323_));
 AOI211_X2 _27338_ (.A(_10900_),
    .B(_05412_),
    .C1(_04605_),
    .C2(_04610_),
    .ZN(_09260_));
 AND2_X1 _27339_ (.A1(_10904_),
    .A2(_09260_),
    .ZN(_09261_));
 BUF_X4 _27340_ (.A(_09261_),
    .Z(_09262_));
 BUF_X4 _27341_ (.A(_09262_),
    .Z(_09263_));
 MUX2_X1 _27342_ (.A(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .B(_06223_),
    .S(_09263_),
    .Z(_02324_));
 MUX2_X1 _27343_ (.A(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .B(_06236_),
    .S(_09263_),
    .Z(_02325_));
 BUF_X4 _27344_ (.A(_09260_),
    .Z(_09264_));
 NAND2_X2 _27345_ (.A1(_10904_),
    .A2(_09264_),
    .ZN(_09265_));
 CLKBUF_X3 _27346_ (.A(_09265_),
    .Z(_09266_));
 NAND2_X1 _27347_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .A2(_09266_),
    .ZN(_09267_));
 OAI21_X1 _27348_ (.A(_09267_),
    .B1(_09266_),
    .B2(_05464_),
    .ZN(_02326_));
 NAND2_X1 _27349_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .A2(_09266_),
    .ZN(_09268_));
 OAI21_X1 _27350_ (.A(_09268_),
    .B1(_09266_),
    .B2(_05510_),
    .ZN(_02327_));
 MUX2_X1 _27351_ (.A(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .B(_09178_),
    .S(_09263_),
    .Z(_02328_));
 MUX2_X1 _27352_ (.A(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .B(_09179_),
    .S(_09263_),
    .Z(_02329_));
 MUX2_X1 _27353_ (.A(_04602_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .S(_06246_),
    .Z(_02330_));
 BUF_X4 _27354_ (.A(_09262_),
    .Z(_09269_));
 MUX2_X1 _27355_ (.A(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .B(_09180_),
    .S(_09269_),
    .Z(_02331_));
 MUX2_X1 _27356_ (.A(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .B(_09181_),
    .S(_09269_),
    .Z(_02332_));
 NOR2_X1 _27357_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .A2(_09263_),
    .ZN(_09270_));
 AOI21_X1 _27358_ (.A(_09270_),
    .B1(_09263_),
    .B2(_05688_),
    .ZN(_02333_));
 MUX2_X1 _27359_ (.A(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .B(_09183_),
    .S(_09269_),
    .Z(_02334_));
 MUX2_X1 _27360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .B(_09185_),
    .S(_09269_),
    .Z(_02335_));
 MUX2_X1 _27361_ (.A(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .B(_09186_),
    .S(_09269_),
    .Z(_02336_));
 NOR2_X1 _27362_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .A2(_09263_),
    .ZN(_09271_));
 AOI21_X1 _27363_ (.A(_09271_),
    .B1(_09263_),
    .B2(_05850_),
    .ZN(_02337_));
 MUX2_X1 _27364_ (.A(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .B(_09188_),
    .S(_09269_),
    .Z(_02338_));
 MUX2_X1 _27365_ (.A(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .B(_09189_),
    .S(_09269_),
    .Z(_02339_));
 MUX2_X1 _27366_ (.A(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .B(_09190_),
    .S(_09269_),
    .Z(_02340_));
 MUX2_X1 _27367_ (.A(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .B(_09198_),
    .S(_09236_),
    .Z(_02341_));
 NOR2_X1 _27368_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .A2(_09263_),
    .ZN(_09272_));
 AOI21_X1 _27369_ (.A(_09272_),
    .B1(_09263_),
    .B2(_06016_),
    .ZN(_02342_));
 MUX2_X1 _27370_ (.A(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .B(_09192_),
    .S(_09269_),
    .Z(_02343_));
 MUX2_X1 _27371_ (.A(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .B(_09193_),
    .S(_09269_),
    .Z(_02344_));
 NAND2_X1 _27372_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .A2(_09266_),
    .ZN(_09273_));
 OAI21_X1 _27373_ (.A(_09273_),
    .B1(_09266_),
    .B2(_06138_),
    .ZN(_02345_));
 MUX2_X1 _27374_ (.A(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .B(_09195_),
    .S(_09262_),
    .Z(_02346_));
 MUX2_X1 _27375_ (.A(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .B(_09196_),
    .S(_09262_),
    .Z(_02347_));
 MUX2_X1 _27376_ (.A(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .B(_09197_),
    .S(_09262_),
    .Z(_02348_));
 MUX2_X1 _27377_ (.A(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .B(_09198_),
    .S(_09262_),
    .Z(_02349_));
 NAND2_X1 _27378_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A2(_09265_),
    .ZN(_09274_));
 OAI21_X1 _27379_ (.A(_09274_),
    .B1(_09266_),
    .B2(_04908_),
    .ZN(_02350_));
 NAND2_X1 _27380_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A2(_09265_),
    .ZN(_09275_));
 OAI21_X4 _27381_ (.A(_09275_),
    .B1(_04978_),
    .B2(_09266_),
    .ZN(_02351_));
 NAND2_X1 _27382_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A2(_09249_),
    .ZN(_09276_));
 OAI21_X1 _27383_ (.A(_09276_),
    .B1(_09251_),
    .B2(_04908_),
    .ZN(_02352_));
 MUX2_X1 _27384_ (.A(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .B(net419),
    .S(_09262_),
    .Z(_02353_));
 MUX2_X1 _27385_ (.A(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .B(net331),
    .S(_09262_),
    .Z(_02354_));
 MUX2_X1 _27386_ (.A(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .B(net408),
    .S(_09262_),
    .Z(_02355_));
 NAND2_X1 _27387_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A2(_09265_),
    .ZN(_09277_));
 OAI21_X4 _27388_ (.A(_09277_),
    .B1(_05148_),
    .B2(_09266_),
    .ZN(_02356_));
 MUX2_X1 _27389_ (.A(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .B(net392),
    .S(_09262_),
    .Z(_02357_));
 NAND2_X1 _27390_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A2(_09265_),
    .ZN(_09278_));
 OAI21_X4 _27391_ (.A(_09278_),
    .B1(_05260_),
    .B2(_09266_),
    .ZN(_02358_));
 AND2_X1 _27392_ (.A1(_06245_),
    .A2(_09260_),
    .ZN(_09279_));
 BUF_X4 _27393_ (.A(_09279_),
    .Z(_09280_));
 BUF_X4 _27394_ (.A(_09280_),
    .Z(_09281_));
 MUX2_X1 _27395_ (.A(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .B(_06223_),
    .S(_09281_),
    .Z(_02359_));
 MUX2_X1 _27396_ (.A(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .B(_06236_),
    .S(_09281_),
    .Z(_02360_));
 NAND2_X2 _27397_ (.A1(_06245_),
    .A2(_09264_),
    .ZN(_09282_));
 CLKBUF_X3 _27398_ (.A(_09282_),
    .Z(_09283_));
 NAND2_X1 _27399_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .A2(_09283_),
    .ZN(_09284_));
 OAI21_X1 _27400_ (.A(_09284_),
    .B1(_09283_),
    .B2(_05464_),
    .ZN(_02361_));
 NAND2_X1 _27401_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .A2(_09283_),
    .ZN(_09285_));
 OAI21_X1 _27402_ (.A(_09285_),
    .B1(_09283_),
    .B2(_05510_),
    .ZN(_02362_));
 NAND2_X1 _27403_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A2(_09249_),
    .ZN(_09286_));
 OAI21_X4 _27404_ (.A(_09286_),
    .B1(_04978_),
    .B2(_09249_),
    .ZN(_02363_));
 MUX2_X1 _27405_ (.A(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .B(_09178_),
    .S(_09281_),
    .Z(_02364_));
 MUX2_X1 _27406_ (.A(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .B(_09179_),
    .S(_09281_),
    .Z(_02365_));
 BUF_X4 _27407_ (.A(_09280_),
    .Z(_09287_));
 MUX2_X1 _27408_ (.A(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .B(_09180_),
    .S(_09287_),
    .Z(_02366_));
 MUX2_X1 _27409_ (.A(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .B(_09181_),
    .S(_09287_),
    .Z(_02367_));
 NOR2_X1 _27410_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .A2(_09281_),
    .ZN(_09288_));
 AOI21_X1 _27411_ (.A(_09288_),
    .B1(_09281_),
    .B2(_05688_),
    .ZN(_02368_));
 MUX2_X1 _27412_ (.A(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .B(_09183_),
    .S(_09287_),
    .Z(_02369_));
 MUX2_X1 _27413_ (.A(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .B(_09185_),
    .S(_09287_),
    .Z(_02370_));
 MUX2_X1 _27414_ (.A(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .B(_09186_),
    .S(_09287_),
    .Z(_02371_));
 NOR2_X1 _27415_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .A2(_09281_),
    .ZN(_09289_));
 AOI21_X1 _27416_ (.A(_09289_),
    .B1(_09281_),
    .B2(_05850_),
    .ZN(_02372_));
 MUX2_X1 _27417_ (.A(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .B(_09188_),
    .S(_09287_),
    .Z(_02373_));
 MUX2_X1 _27418_ (.A(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B(_09201_),
    .S(_09236_),
    .Z(_02374_));
 MUX2_X1 _27419_ (.A(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .B(_09189_),
    .S(_09287_),
    .Z(_02375_));
 MUX2_X1 _27420_ (.A(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .B(_09190_),
    .S(_09287_),
    .Z(_02376_));
 NOR2_X1 _27421_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .A2(_09281_),
    .ZN(_09290_));
 AOI21_X1 _27422_ (.A(_09290_),
    .B1(_09281_),
    .B2(_06016_),
    .ZN(_02377_));
 MUX2_X1 _27423_ (.A(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .B(_09192_),
    .S(_09287_),
    .Z(_02378_));
 MUX2_X1 _27424_ (.A(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .B(_09193_),
    .S(_09287_),
    .Z(_02379_));
 NAND2_X1 _27425_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .A2(_09283_),
    .ZN(_09291_));
 CLKBUF_X3 _27426_ (.A(_06137_),
    .Z(_09292_));
 OAI21_X1 _27427_ (.A(_09291_),
    .B1(_09283_),
    .B2(_09292_),
    .ZN(_02380_));
 MUX2_X1 _27428_ (.A(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .B(_09195_),
    .S(_09280_),
    .Z(_02381_));
 MUX2_X1 _27429_ (.A(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .B(_09196_),
    .S(_09280_),
    .Z(_02382_));
 MUX2_X1 _27430_ (.A(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .B(_09197_),
    .S(_09280_),
    .Z(_02383_));
 MUX2_X1 _27431_ (.A(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .B(_09198_),
    .S(_09280_),
    .Z(_02384_));
 BUF_X4 _27432_ (.A(_04849_),
    .Z(_09293_));
 MUX2_X1 _27433_ (.A(net332),
    .B(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .S(_06246_),
    .Z(_02385_));
 NAND2_X1 _27434_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .A2(_09282_),
    .ZN(_09294_));
 BUF_X8 _27435_ (.A(_04907_),
    .Z(_09295_));
 OAI21_X1 _27436_ (.A(_09294_),
    .B1(_09283_),
    .B2(_09295_),
    .ZN(_02386_));
 NAND2_X1 _27437_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .A2(_09282_),
    .ZN(_09296_));
 BUF_X8 _27438_ (.A(_04977_),
    .Z(_09297_));
 OAI21_X1 _27439_ (.A(_09296_),
    .B1(_09283_),
    .B2(_09297_),
    .ZN(_02387_));
 MUX2_X1 _27440_ (.A(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .B(_09201_),
    .S(_09280_),
    .Z(_02388_));
 MUX2_X1 _27441_ (.A(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .B(_09202_),
    .S(_09280_),
    .Z(_02389_));
 MUX2_X1 _27442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .B(net408),
    .S(_09280_),
    .Z(_02390_));
 NAND2_X1 _27443_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .A2(_09282_),
    .ZN(_09298_));
 OAI21_X4 _27444_ (.A(_09298_),
    .B1(_05148_),
    .B2(_09283_),
    .ZN(_02391_));
 MUX2_X1 _27445_ (.A(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .B(_06208_),
    .S(_09280_),
    .Z(_02392_));
 NAND2_X1 _27446_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A2(_09282_),
    .ZN(_09299_));
 OAI21_X4 _27447_ (.A(_09299_),
    .B1(_05260_),
    .B2(_09283_),
    .ZN(_02393_));
 NOR2_X4 _27448_ (.A1(_10903_),
    .A2(_05373_),
    .ZN(_09300_));
 AND2_X1 _27449_ (.A1(_09264_),
    .A2(_09300_),
    .ZN(_09301_));
 BUF_X4 _27450_ (.A(_09301_),
    .Z(_09302_));
 BUF_X4 _27451_ (.A(_09302_),
    .Z(_09303_));
 MUX2_X1 _27452_ (.A(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .B(_06223_),
    .S(_09303_),
    .Z(_02394_));
 MUX2_X1 _27453_ (.A(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .B(_06236_),
    .S(_09303_),
    .Z(_02395_));
 MUX2_X1 _27454_ (.A(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .B(_05411_),
    .S(_09236_),
    .Z(_02396_));
 NAND2_X2 _27455_ (.A1(_09264_),
    .A2(_09300_),
    .ZN(_09304_));
 BUF_X4 _27456_ (.A(_09304_),
    .Z(_09305_));
 NAND2_X1 _27457_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .A2(_09305_),
    .ZN(_09306_));
 CLKBUF_X3 _27458_ (.A(_05463_),
    .Z(_09307_));
 OAI21_X1 _27459_ (.A(_09306_),
    .B1(_09305_),
    .B2(_09307_),
    .ZN(_02397_));
 NAND2_X1 _27460_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .A2(_09305_),
    .ZN(_09308_));
 CLKBUF_X3 _27461_ (.A(_05509_),
    .Z(_09309_));
 OAI21_X1 _27462_ (.A(_09308_),
    .B1(_09305_),
    .B2(_09309_),
    .ZN(_02398_));
 MUX2_X1 _27463_ (.A(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .B(_09178_),
    .S(_09303_),
    .Z(_02399_));
 MUX2_X1 _27464_ (.A(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .B(_09179_),
    .S(_09303_),
    .Z(_02400_));
 BUF_X4 _27465_ (.A(_09302_),
    .Z(_09310_));
 MUX2_X1 _27466_ (.A(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .B(_09180_),
    .S(_09310_),
    .Z(_02401_));
 MUX2_X1 _27467_ (.A(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .B(_09181_),
    .S(_09310_),
    .Z(_02402_));
 NOR2_X1 _27468_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .A2(_09303_),
    .ZN(_09311_));
 AOI21_X1 _27469_ (.A(_09311_),
    .B1(_09303_),
    .B2(_05688_),
    .ZN(_02403_));
 MUX2_X1 _27470_ (.A(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .B(_09183_),
    .S(_09310_),
    .Z(_02404_));
 MUX2_X1 _27471_ (.A(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .B(_09185_),
    .S(_09310_),
    .Z(_02405_));
 MUX2_X1 _27472_ (.A(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .B(_09186_),
    .S(_09310_),
    .Z(_02406_));
 NAND2_X1 _27473_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A2(_09249_),
    .ZN(_09312_));
 BUF_X8 _27474_ (.A(_05147_),
    .Z(_09313_));
 OAI21_X4 _27475_ (.A(_09312_),
    .B1(net444),
    .B2(_09251_),
    .ZN(_02407_));
 NAND2_X1 _27476_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .A2(_09249_),
    .ZN(_09314_));
 OAI21_X1 _27477_ (.A(_09314_),
    .B1(_09249_),
    .B2(_09307_),
    .ZN(_02408_));
 NOR2_X1 _27478_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .A2(_09303_),
    .ZN(_09315_));
 CLKBUF_X3 _27479_ (.A(_05849_),
    .Z(_09316_));
 AOI21_X1 _27480_ (.A(_09315_),
    .B1(_09303_),
    .B2(_09316_),
    .ZN(_02409_));
 MUX2_X1 _27481_ (.A(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .B(_09188_),
    .S(_09310_),
    .Z(_02410_));
 MUX2_X1 _27482_ (.A(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .B(_09189_),
    .S(_09310_),
    .Z(_02411_));
 MUX2_X1 _27483_ (.A(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .B(_09190_),
    .S(_09310_),
    .Z(_02412_));
 NOR2_X1 _27484_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .A2(_09303_),
    .ZN(_09317_));
 CLKBUF_X3 _27485_ (.A(_06015_),
    .Z(_09318_));
 AOI21_X1 _27486_ (.A(_09317_),
    .B1(_09303_),
    .B2(_09318_),
    .ZN(_02413_));
 MUX2_X1 _27487_ (.A(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .B(_09192_),
    .S(_09310_),
    .Z(_02414_));
 MUX2_X1 _27488_ (.A(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .B(_09193_),
    .S(_09310_),
    .Z(_02415_));
 NAND2_X1 _27489_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .A2(_09305_),
    .ZN(_09319_));
 OAI21_X1 _27490_ (.A(_09319_),
    .B1(_09305_),
    .B2(_09292_),
    .ZN(_02416_));
 MUX2_X1 _27491_ (.A(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .B(_09195_),
    .S(_09302_),
    .Z(_02417_));
 MUX2_X1 _27492_ (.A(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .B(_09196_),
    .S(_09302_),
    .Z(_02418_));
 MUX2_X1 _27493_ (.A(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .B(_06208_),
    .S(_09236_),
    .Z(_02419_));
 MUX2_X1 _27494_ (.A(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .B(_09197_),
    .S(_09302_),
    .Z(_02420_));
 MUX2_X1 _27495_ (.A(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .B(_09198_),
    .S(_09302_),
    .Z(_02421_));
 NAND2_X1 _27496_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A2(_09304_),
    .ZN(_09320_));
 OAI21_X1 _27497_ (.A(_09320_),
    .B1(_09305_),
    .B2(net412),
    .ZN(_02422_));
 NAND2_X1 _27498_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .A2(_09304_),
    .ZN(_09321_));
 OAI21_X1 _27499_ (.A(_09321_),
    .B1(_09305_),
    .B2(_09297_),
    .ZN(_02423_));
 MUX2_X1 _27500_ (.A(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .B(_09201_),
    .S(_09302_),
    .Z(_02424_));
 MUX2_X1 _27501_ (.A(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .B(net331),
    .S(_09302_),
    .Z(_02425_));
 MUX2_X1 _27502_ (.A(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .B(_05411_),
    .S(_09302_),
    .Z(_02426_));
 NAND2_X1 _27503_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .A2(_09304_),
    .ZN(_09322_));
 OAI21_X4 _27504_ (.A(_09322_),
    .B1(_09313_),
    .B2(_09305_),
    .ZN(_02427_));
 MUX2_X1 _27505_ (.A(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .B(_06208_),
    .S(_09302_),
    .Z(_02428_));
 NAND2_X1 _27506_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A2(_09304_),
    .ZN(_09323_));
 BUF_X8 _27507_ (.A(_05259_),
    .Z(_09324_));
 OAI21_X2 _27508_ (.A(_09323_),
    .B1(_09305_),
    .B2(_09324_),
    .ZN(_02429_));
 NAND2_X1 _27509_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A2(_09249_),
    .ZN(_09325_));
 OAI21_X2 _27510_ (.A(_09325_),
    .B1(net422),
    .B2(_09251_),
    .ZN(_02430_));
 AND2_X1 _27511_ (.A1(_04852_),
    .A2(_09260_),
    .ZN(_09326_));
 BUF_X4 _27512_ (.A(_09326_),
    .Z(_09327_));
 BUF_X4 _27513_ (.A(_09327_),
    .Z(_09328_));
 MUX2_X1 _27514_ (.A(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .B(_06223_),
    .S(_09328_),
    .Z(_02431_));
 MUX2_X1 _27515_ (.A(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .B(_06236_),
    .S(_09328_),
    .Z(_02432_));
 NAND2_X2 _27516_ (.A1(_04852_),
    .A2(_09264_),
    .ZN(_09329_));
 CLKBUF_X3 _27517_ (.A(_09329_),
    .Z(_09330_));
 NAND2_X1 _27518_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .A2(_09330_),
    .ZN(_09331_));
 OAI21_X1 _27519_ (.A(_09331_),
    .B1(_09330_),
    .B2(_09307_),
    .ZN(_02433_));
 NAND2_X1 _27520_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .A2(_09330_),
    .ZN(_09332_));
 OAI21_X1 _27521_ (.A(_09332_),
    .B1(_09330_),
    .B2(_09309_),
    .ZN(_02434_));
 MUX2_X1 _27522_ (.A(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .B(_09178_),
    .S(_09328_),
    .Z(_02435_));
 MUX2_X1 _27523_ (.A(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .B(_09179_),
    .S(_09328_),
    .Z(_02436_));
 BUF_X4 _27524_ (.A(_09327_),
    .Z(_09333_));
 MUX2_X1 _27525_ (.A(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .B(_09180_),
    .S(_09333_),
    .Z(_02437_));
 MUX2_X1 _27526_ (.A(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .B(_09181_),
    .S(_09333_),
    .Z(_02438_));
 NOR2_X1 _27527_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .A2(_09328_),
    .ZN(_09334_));
 AOI21_X1 _27528_ (.A(_09334_),
    .B1(_09328_),
    .B2(_05688_),
    .ZN(_02439_));
 MUX2_X1 _27529_ (.A(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .B(_09183_),
    .S(_09333_),
    .Z(_02440_));
 AND2_X1 _27530_ (.A1(_05805_),
    .A2(_09300_),
    .ZN(_09335_));
 BUF_X4 _27531_ (.A(_09335_),
    .Z(_09336_));
 MUX2_X1 _27532_ (.A(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .B(_06223_),
    .S(_09336_),
    .Z(_02441_));
 MUX2_X1 _27533_ (.A(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .B(_09185_),
    .S(_09333_),
    .Z(_02442_));
 MUX2_X1 _27534_ (.A(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .B(_09186_),
    .S(_09333_),
    .Z(_02443_));
 NOR2_X1 _27535_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .A2(_09328_),
    .ZN(_09337_));
 AOI21_X1 _27536_ (.A(_09337_),
    .B1(_09328_),
    .B2(_09316_),
    .ZN(_02444_));
 MUX2_X1 _27537_ (.A(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .B(_09188_),
    .S(_09333_),
    .Z(_02445_));
 MUX2_X1 _27538_ (.A(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .B(_09189_),
    .S(_09333_),
    .Z(_02446_));
 MUX2_X1 _27539_ (.A(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .B(_09190_),
    .S(_09333_),
    .Z(_02447_));
 NOR2_X1 _27540_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .A2(_09328_),
    .ZN(_09338_));
 AOI21_X1 _27541_ (.A(_09338_),
    .B1(_09328_),
    .B2(_09318_),
    .ZN(_02448_));
 MUX2_X1 _27542_ (.A(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .B(_09192_),
    .S(_09333_),
    .Z(_02449_));
 MUX2_X1 _27543_ (.A(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .B(_09193_),
    .S(_09333_),
    .Z(_02450_));
 NAND2_X1 _27544_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .A2(_09330_),
    .ZN(_09339_));
 OAI21_X1 _27545_ (.A(_09339_),
    .B1(_09330_),
    .B2(_09292_),
    .ZN(_02451_));
 MUX2_X1 _27546_ (.A(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .B(_06236_),
    .S(_09336_),
    .Z(_02452_));
 MUX2_X1 _27547_ (.A(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .B(_09195_),
    .S(_09327_),
    .Z(_02453_));
 MUX2_X1 _27548_ (.A(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .B(_09196_),
    .S(_09327_),
    .Z(_02454_));
 MUX2_X1 _27549_ (.A(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .B(_09197_),
    .S(_09327_),
    .Z(_02455_));
 MUX2_X1 _27550_ (.A(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .B(_09198_),
    .S(_09327_),
    .Z(_02456_));
 NAND2_X1 _27551_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .A2(_09329_),
    .ZN(_09340_));
 OAI21_X1 _27552_ (.A(_09340_),
    .B1(_09330_),
    .B2(_09295_),
    .ZN(_02457_));
 NAND2_X1 _27553_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .A2(_09329_),
    .ZN(_09341_));
 OAI21_X1 _27554_ (.A(_09341_),
    .B1(_09330_),
    .B2(_09297_),
    .ZN(_02458_));
 MUX2_X1 _27555_ (.A(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .B(net419),
    .S(_09327_),
    .Z(_02459_));
 MUX2_X1 _27556_ (.A(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .B(net331),
    .S(_09327_),
    .Z(_02460_));
 MUX2_X1 _27557_ (.A(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .B(_05411_),
    .S(_09327_),
    .Z(_02461_));
 NAND2_X1 _27558_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .A2(_09329_),
    .ZN(_09342_));
 OAI21_X4 _27559_ (.A(_09342_),
    .B1(net444),
    .B2(_09330_),
    .ZN(_02462_));
 NAND2_X4 _27560_ (.A1(_04854_),
    .A2(_09300_),
    .ZN(_09343_));
 CLKBUF_X3 _27561_ (.A(_09343_),
    .Z(_09344_));
 NAND2_X1 _27562_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A2(_09344_),
    .ZN(_09345_));
 OAI21_X1 _27563_ (.A(_09345_),
    .B1(_09344_),
    .B2(_09307_),
    .ZN(_02463_));
 MUX2_X1 _27564_ (.A(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .B(net392),
    .S(_09327_),
    .Z(_02464_));
 NAND2_X1 _27565_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .A2(_09329_),
    .ZN(_09346_));
 OAI21_X2 _27566_ (.A(_09346_),
    .B1(_09330_),
    .B2(_09324_),
    .ZN(_02465_));
 NAND2_X4 _27567_ (.A1(_10904_),
    .A2(_04613_),
    .ZN(_09347_));
 BUF_X4 _27568_ (.A(_09347_),
    .Z(_09348_));
 MUX2_X1 _27569_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .S(_09348_),
    .Z(_02466_));
 MUX2_X1 _27570_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .S(_09348_),
    .Z(_02467_));
 BUF_X4 _27571_ (.A(_09347_),
    .Z(_09349_));
 NAND2_X1 _27572_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .A2(_09349_),
    .ZN(_09350_));
 BUF_X4 _27573_ (.A(_09347_),
    .Z(_09351_));
 OAI21_X1 _27574_ (.A(_09350_),
    .B1(_09351_),
    .B2(_09307_),
    .ZN(_02468_));
 NAND2_X1 _27575_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .A2(_09349_),
    .ZN(_09352_));
 OAI21_X1 _27576_ (.A(_09352_),
    .B1(_09351_),
    .B2(_09309_),
    .ZN(_02469_));
 MUX2_X1 _27577_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .S(_09348_),
    .Z(_02470_));
 MUX2_X1 _27578_ (.A(_05580_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .S(_09348_),
    .Z(_02471_));
 MUX2_X1 _27579_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .S(_09348_),
    .Z(_02472_));
 MUX2_X1 _27580_ (.A(_05653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .S(_09348_),
    .Z(_02473_));
 NAND2_X1 _27581_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .A2(_09344_),
    .ZN(_09353_));
 OAI21_X1 _27582_ (.A(_09353_),
    .B1(_09344_),
    .B2(_09309_),
    .ZN(_02474_));
 NAND2_X1 _27583_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .A2(_09349_),
    .ZN(_09354_));
 OAI21_X1 _27584_ (.A(_09354_),
    .B1(_09351_),
    .B2(_06222_),
    .ZN(_02475_));
 MUX2_X1 _27585_ (.A(_05721_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .S(_09348_),
    .Z(_02476_));
 MUX2_X1 _27586_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .S(_09348_),
    .Z(_02477_));
 MUX2_X1 _27587_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .S(_09348_),
    .Z(_02478_));
 NAND2_X1 _27588_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .A2(_09349_),
    .ZN(_09355_));
 OAI21_X1 _27589_ (.A(_09355_),
    .B1(_09351_),
    .B2(_06231_),
    .ZN(_02479_));
 MUX2_X1 _27590_ (.A(_05890_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .S(_09348_),
    .Z(_02480_));
 BUF_X4 _27591_ (.A(_09347_),
    .Z(_09356_));
 MUX2_X1 _27592_ (.A(_05928_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .S(_09356_),
    .Z(_02481_));
 MUX2_X1 _27593_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .S(_09356_),
    .Z(_02482_));
 NAND2_X1 _27594_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .A2(_09349_),
    .ZN(_09357_));
 OAI21_X1 _27595_ (.A(_09357_),
    .B1(_09351_),
    .B2(_06234_),
    .ZN(_02483_));
 MUX2_X1 _27596_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .S(_09356_),
    .Z(_02484_));
 MUX2_X1 _27597_ (.A(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .B(_09178_),
    .S(_09336_),
    .Z(_02485_));
 MUX2_X1 _27598_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .S(_09356_),
    .Z(_02486_));
 NAND2_X1 _27599_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .A2(_09349_),
    .ZN(_09358_));
 OAI21_X1 _27600_ (.A(_09358_),
    .B1(_09351_),
    .B2(_09292_),
    .ZN(_02487_));
 MUX2_X1 _27601_ (.A(_06174_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .S(_09356_),
    .Z(_02488_));
 MUX2_X1 _27602_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .S(_09356_),
    .Z(_02489_));
 BUF_X2 _27603_ (.A(_04601_),
    .Z(_09359_));
 MUX2_X1 _27604_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .S(_09356_),
    .Z(_02490_));
 MUX2_X1 _27605_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .S(_09356_),
    .Z(_02491_));
 NAND2_X1 _27606_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A2(_09349_),
    .ZN(_09360_));
 OAI21_X1 _27607_ (.A(_09360_),
    .B1(_09351_),
    .B2(_09295_),
    .ZN(_02492_));
 NAND2_X1 _27608_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A2(_09349_),
    .ZN(_09361_));
 OAI21_X1 _27609_ (.A(_09361_),
    .B1(_09351_),
    .B2(_09297_),
    .ZN(_02493_));
 MUX2_X1 _27610_ (.A(_05037_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .S(_09356_),
    .Z(_02494_));
 MUX2_X1 _27611_ (.A(_09293_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .S(_09356_),
    .Z(_02495_));
 MUX2_X1 _27612_ (.A(_05580_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .S(_09343_),
    .Z(_02496_));
 MUX2_X1 _27613_ (.A(net409),
    .B(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .S(_09347_),
    .Z(_02497_));
 NAND2_X1 _27614_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A2(_09349_),
    .ZN(_09362_));
 OAI21_X1 _27615_ (.A(_09362_),
    .B1(_09351_),
    .B2(_09313_),
    .ZN(_02498_));
 MUX2_X1 _27616_ (.A(_05211_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .S(_09347_),
    .Z(_02499_));
 NAND2_X1 _27617_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A2(_09349_),
    .ZN(_09363_));
 OAI21_X4 _27618_ (.A(_09363_),
    .B1(_09324_),
    .B2(_09351_),
    .ZN(_02500_));
 NAND2_X4 _27619_ (.A1(_04613_),
    .A2(_06245_),
    .ZN(_09364_));
 BUF_X4 _27620_ (.A(_09364_),
    .Z(_09365_));
 MUX2_X1 _27621_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .S(_09365_),
    .Z(_02501_));
 MUX2_X1 _27622_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .S(_09365_),
    .Z(_02502_));
 BUF_X4 _27623_ (.A(_09364_),
    .Z(_09366_));
 NAND2_X1 _27624_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .A2(_09366_),
    .ZN(_09367_));
 BUF_X4 _27625_ (.A(_09364_),
    .Z(_09368_));
 OAI21_X1 _27626_ (.A(_09367_),
    .B1(_09368_),
    .B2(_09307_),
    .ZN(_02503_));
 NAND2_X1 _27627_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .A2(_09366_),
    .ZN(_09369_));
 OAI21_X1 _27628_ (.A(_09369_),
    .B1(_09368_),
    .B2(_09309_),
    .ZN(_02504_));
 MUX2_X1 _27629_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .S(_09365_),
    .Z(_02505_));
 BUF_X2 _27630_ (.A(_05579_),
    .Z(_09370_));
 MUX2_X1 _27631_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .S(_09365_),
    .Z(_02506_));
 MUX2_X1 _27632_ (.A(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .B(_09180_),
    .S(_09336_),
    .Z(_02507_));
 MUX2_X1 _27633_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .S(_09365_),
    .Z(_02508_));
 MUX2_X1 _27634_ (.A(_05653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .S(_09365_),
    .Z(_02509_));
 NAND2_X1 _27635_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .A2(_09366_),
    .ZN(_09371_));
 OAI21_X1 _27636_ (.A(_09371_),
    .B1(_09368_),
    .B2(_06222_),
    .ZN(_02510_));
 BUF_X2 _27637_ (.A(_05720_),
    .Z(_09372_));
 MUX2_X1 _27638_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .S(_09365_),
    .Z(_02511_));
 MUX2_X1 _27639_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .S(_09365_),
    .Z(_02512_));
 MUX2_X1 _27640_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .S(_09365_),
    .Z(_02513_));
 NAND2_X1 _27641_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .A2(_09366_),
    .ZN(_09373_));
 OAI21_X1 _27642_ (.A(_09373_),
    .B1(_09368_),
    .B2(_06231_),
    .ZN(_02514_));
 BUF_X2 _27643_ (.A(_05889_),
    .Z(_09374_));
 MUX2_X1 _27644_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .S(_09365_),
    .Z(_02515_));
 BUF_X2 _27645_ (.A(_05927_),
    .Z(_09375_));
 BUF_X4 _27646_ (.A(_09364_),
    .Z(_09376_));
 MUX2_X1 _27647_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .S(_09376_),
    .Z(_02516_));
 MUX2_X1 _27648_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .S(_09376_),
    .Z(_02517_));
 BUF_X2 _27649_ (.A(_05652_),
    .Z(_09377_));
 MUX2_X1 _27650_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .S(_09343_),
    .Z(_02518_));
 NAND2_X1 _27651_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .A2(_09249_),
    .ZN(_09378_));
 OAI21_X1 _27652_ (.A(_09378_),
    .B1(_09249_),
    .B2(_09309_),
    .ZN(_02519_));
 NAND2_X1 _27653_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .A2(_09366_),
    .ZN(_09379_));
 OAI21_X1 _27654_ (.A(_09379_),
    .B1(_09368_),
    .B2(_06234_),
    .ZN(_02520_));
 MUX2_X1 _27655_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .S(_09376_),
    .Z(_02521_));
 MUX2_X1 _27656_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .S(_09376_),
    .Z(_02522_));
 NAND2_X1 _27657_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .A2(_09366_),
    .ZN(_09380_));
 OAI21_X1 _27658_ (.A(_09380_),
    .B1(_09368_),
    .B2(_09292_),
    .ZN(_02523_));
 MUX2_X1 _27659_ (.A(net405),
    .B(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .S(_09376_),
    .Z(_02524_));
 MUX2_X1 _27660_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .S(_09376_),
    .Z(_02525_));
 MUX2_X1 _27661_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .S(_09376_),
    .Z(_02526_));
 MUX2_X1 _27662_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .S(_09376_),
    .Z(_02527_));
 NAND2_X1 _27663_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .A2(_09366_),
    .ZN(_09381_));
 OAI21_X1 _27664_ (.A(_09381_),
    .B1(_09368_),
    .B2(net412),
    .ZN(_02528_));
 NAND2_X1 _27665_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .A2(_09366_),
    .ZN(_09382_));
 OAI21_X1 _27666_ (.A(_09382_),
    .B1(_09368_),
    .B2(_09297_),
    .ZN(_02529_));
 NOR2_X1 _27667_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A2(_09336_),
    .ZN(_09383_));
 CLKBUF_X3 _27668_ (.A(_05687_),
    .Z(_09384_));
 AOI21_X1 _27669_ (.A(_09383_),
    .B1(_09336_),
    .B2(_09384_),
    .ZN(_02530_));
 MUX2_X1 _27670_ (.A(net418),
    .B(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .S(_09376_),
    .Z(_02531_));
 MUX2_X1 _27671_ (.A(net332),
    .B(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .S(_09376_),
    .Z(_02532_));
 MUX2_X1 _27672_ (.A(net409),
    .B(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .S(_09364_),
    .Z(_02533_));
 NAND2_X1 _27673_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .A2(_09366_),
    .ZN(_09385_));
 OAI21_X4 _27674_ (.A(_09385_),
    .B1(_09313_),
    .B2(_09368_),
    .ZN(_02534_));
 MUX2_X1 _27675_ (.A(net400),
    .B(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .S(_09364_),
    .Z(_02535_));
 NAND2_X1 _27676_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .A2(_09366_),
    .ZN(_09386_));
 OAI21_X2 _27677_ (.A(_09386_),
    .B1(_09368_),
    .B2(_09324_),
    .ZN(_02536_));
 NAND2_X4 _27678_ (.A1(_04613_),
    .A2(_09300_),
    .ZN(_09387_));
 BUF_X4 _27679_ (.A(_09387_),
    .Z(_09388_));
 MUX2_X1 _27680_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S(_09388_),
    .Z(_02537_));
 MUX2_X1 _27681_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .S(_09388_),
    .Z(_02538_));
 BUF_X4 _27682_ (.A(_09387_),
    .Z(_09389_));
 NAND2_X1 _27683_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .A2(_09389_),
    .ZN(_09390_));
 BUF_X4 _27684_ (.A(_09387_),
    .Z(_09391_));
 OAI21_X1 _27685_ (.A(_09390_),
    .B1(_09391_),
    .B2(_09307_),
    .ZN(_02539_));
 NAND2_X1 _27686_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .A2(_09389_),
    .ZN(_09392_));
 OAI21_X1 _27687_ (.A(_09392_),
    .B1(_09391_),
    .B2(_09309_),
    .ZN(_02540_));
 MUX2_X1 _27688_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .S(_09343_),
    .Z(_02541_));
 MUX2_X1 _27689_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .S(_09388_),
    .Z(_02542_));
 MUX2_X1 _27690_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S(_09388_),
    .Z(_02543_));
 MUX2_X1 _27691_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S(_09388_),
    .Z(_02544_));
 MUX2_X1 _27692_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S(_09388_),
    .Z(_02545_));
 NAND2_X1 _27693_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .A2(_09389_),
    .ZN(_09393_));
 OAI21_X1 _27694_ (.A(_09393_),
    .B1(_09391_),
    .B2(_06222_),
    .ZN(_02546_));
 MUX2_X1 _27695_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S(_09388_),
    .Z(_02547_));
 MUX2_X1 _27696_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S(_09388_),
    .Z(_02548_));
 MUX2_X1 _27697_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(_09388_),
    .Z(_02549_));
 NAND2_X1 _27698_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .A2(_09389_),
    .ZN(_09394_));
 OAI21_X1 _27699_ (.A(_09394_),
    .B1(_09391_),
    .B2(_06231_),
    .ZN(_02550_));
 MUX2_X1 _27700_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .S(_09388_),
    .Z(_02551_));
 BUF_X4 _27701_ (.A(_09335_),
    .Z(_09395_));
 MUX2_X1 _27702_ (.A(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .B(_09185_),
    .S(_09395_),
    .Z(_02552_));
 BUF_X4 _27703_ (.A(_09387_),
    .Z(_09396_));
 MUX2_X1 _27704_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .S(_09396_),
    .Z(_02553_));
 MUX2_X1 _27705_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .S(_09396_),
    .Z(_02554_));
 NAND2_X1 _27706_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .A2(_09389_),
    .ZN(_09397_));
 OAI21_X1 _27707_ (.A(_09397_),
    .B1(_09391_),
    .B2(_06234_),
    .ZN(_02555_));
 MUX2_X1 _27708_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .S(_09396_),
    .Z(_02556_));
 MUX2_X1 _27709_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .S(_09396_),
    .Z(_02557_));
 NAND2_X1 _27710_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .A2(_09389_),
    .ZN(_09398_));
 OAI21_X1 _27711_ (.A(_09398_),
    .B1(_09391_),
    .B2(_09292_),
    .ZN(_02558_));
 MUX2_X1 _27712_ (.A(_06174_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .S(_09396_),
    .Z(_02559_));
 MUX2_X1 _27713_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .S(_09396_),
    .Z(_02560_));
 MUX2_X1 _27714_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .S(_09396_),
    .Z(_02561_));
 MUX2_X1 _27715_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .S(_09396_),
    .Z(_02562_));
 MUX2_X1 _27716_ (.A(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .B(_09186_),
    .S(_09395_),
    .Z(_02563_));
 NAND2_X1 _27717_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A2(_09389_),
    .ZN(_09399_));
 OAI21_X1 _27718_ (.A(_09399_),
    .B1(_09391_),
    .B2(_09295_),
    .ZN(_02564_));
 NAND2_X1 _27719_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .A2(_09389_),
    .ZN(_09400_));
 OAI21_X1 _27720_ (.A(_09400_),
    .B1(_09391_),
    .B2(_09297_),
    .ZN(_02565_));
 MUX2_X1 _27721_ (.A(net418),
    .B(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .S(_09396_),
    .Z(_02566_));
 MUX2_X1 _27722_ (.A(_09293_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .S(_09396_),
    .Z(_02567_));
 MUX2_X1 _27723_ (.A(_05094_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .S(_09387_),
    .Z(_02568_));
 NAND2_X1 _27724_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .A2(_09389_),
    .ZN(_09401_));
 OAI21_X1 _27725_ (.A(_09401_),
    .B1(_09391_),
    .B2(_09313_),
    .ZN(_02569_));
 MUX2_X1 _27726_ (.A(net400),
    .B(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .S(_09387_),
    .Z(_02570_));
 NAND2_X1 _27727_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A2(_09389_),
    .ZN(_09402_));
 OAI21_X2 _27728_ (.A(_09402_),
    .B1(net422),
    .B2(_09391_),
    .ZN(_02571_));
 NAND2_X4 _27729_ (.A1(_04613_),
    .A2(_04852_),
    .ZN(_09403_));
 BUF_X4 _27730_ (.A(_09403_),
    .Z(_09404_));
 MUX2_X1 _27731_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(_09404_),
    .Z(_02572_));
 MUX2_X1 _27732_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S(_09404_),
    .Z(_02573_));
 NOR2_X1 _27733_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A2(_09336_),
    .ZN(_09405_));
 AOI21_X1 _27734_ (.A(_09405_),
    .B1(_09336_),
    .B2(_09316_),
    .ZN(_02574_));
 BUF_X4 _27735_ (.A(_09403_),
    .Z(_09406_));
 NAND2_X1 _27736_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .A2(_09406_),
    .ZN(_09407_));
 BUF_X4 _27737_ (.A(_09403_),
    .Z(_09408_));
 OAI21_X1 _27738_ (.A(_09407_),
    .B1(_09408_),
    .B2(_09307_),
    .ZN(_02575_));
 NAND2_X1 _27739_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .A2(_09406_),
    .ZN(_09409_));
 OAI21_X1 _27740_ (.A(_09409_),
    .B1(_09408_),
    .B2(_09309_),
    .ZN(_02576_));
 MUX2_X1 _27741_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(_09404_),
    .Z(_02577_));
 MUX2_X1 _27742_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(_09404_),
    .Z(_02578_));
 MUX2_X1 _27743_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S(_09404_),
    .Z(_02579_));
 MUX2_X1 _27744_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(_09404_),
    .Z(_02580_));
 NAND2_X1 _27745_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .A2(_09406_),
    .ZN(_09410_));
 OAI21_X1 _27746_ (.A(_09410_),
    .B1(_09408_),
    .B2(_06222_),
    .ZN(_02581_));
 MUX2_X1 _27747_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(_09404_),
    .Z(_02582_));
 MUX2_X1 _27748_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(_09404_),
    .Z(_02583_));
 MUX2_X1 _27749_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(_09404_),
    .Z(_02584_));
 MUX2_X1 _27750_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .S(_09343_),
    .Z(_02585_));
 NAND2_X1 _27751_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .A2(_09406_),
    .ZN(_09411_));
 OAI21_X1 _27752_ (.A(_09411_),
    .B1(_09408_),
    .B2(_06231_),
    .ZN(_02586_));
 MUX2_X1 _27753_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(_09404_),
    .Z(_02587_));
 BUF_X4 _27754_ (.A(_09403_),
    .Z(_09412_));
 MUX2_X1 _27755_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S(_09412_),
    .Z(_02588_));
 MUX2_X1 _27756_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(_09412_),
    .Z(_02589_));
 NAND2_X1 _27757_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .A2(_09406_),
    .ZN(_09413_));
 OAI21_X1 _27758_ (.A(_09413_),
    .B1(_09408_),
    .B2(_06234_),
    .ZN(_02590_));
 MUX2_X1 _27759_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S(_09412_),
    .Z(_02591_));
 MUX2_X1 _27760_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S(_09412_),
    .Z(_02592_));
 NAND2_X1 _27761_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .A2(_09406_),
    .ZN(_09414_));
 OAI21_X1 _27762_ (.A(_09414_),
    .B1(_09408_),
    .B2(_09292_),
    .ZN(_02593_));
 MUX2_X1 _27763_ (.A(net405),
    .B(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S(_09412_),
    .Z(_02594_));
 MUX2_X1 _27764_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S(_09412_),
    .Z(_02595_));
 MUX2_X1 _27765_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .S(_09343_),
    .Z(_02596_));
 MUX2_X1 _27766_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S(_09412_),
    .Z(_02597_));
 MUX2_X1 _27767_ (.A(_04766_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S(_09412_),
    .Z(_02598_));
 NAND2_X1 _27768_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .A2(_09406_),
    .ZN(_09415_));
 OAI21_X1 _27769_ (.A(_09415_),
    .B1(_09408_),
    .B2(_09295_),
    .ZN(_02599_));
 NAND2_X1 _27770_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .A2(_09406_),
    .ZN(_09416_));
 OAI21_X1 _27771_ (.A(_09416_),
    .B1(_09408_),
    .B2(_09297_),
    .ZN(_02600_));
 MUX2_X1 _27772_ (.A(_05037_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(_09412_),
    .Z(_02601_));
 MUX2_X1 _27773_ (.A(net332),
    .B(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S(_09412_),
    .Z(_02602_));
 MUX2_X1 _27774_ (.A(net409),
    .B(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S(_09403_),
    .Z(_02603_));
 NAND2_X1 _27775_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .A2(_09406_),
    .ZN(_09417_));
 OAI21_X4 _27776_ (.A(_09417_),
    .B1(_09313_),
    .B2(_09408_),
    .ZN(_02604_));
 MUX2_X1 _27777_ (.A(_05211_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S(_09403_),
    .Z(_02605_));
 NAND2_X1 _27778_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .A2(_09406_),
    .ZN(_09418_));
 OAI21_X4 _27779_ (.A(_09418_),
    .B1(_09324_),
    .B2(_09408_),
    .ZN(_02606_));
 MUX2_X1 _27780_ (.A(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .B(_09190_),
    .S(_09395_),
    .Z(_02607_));
 BUF_X2 _27781_ (.A(_05371_),
    .Z(_09419_));
 NOR3_X4 _27782_ (.A1(_10394_),
    .A2(_10902_),
    .A3(_04603_),
    .ZN(_09420_));
 AND2_X1 _27783_ (.A1(_05805_),
    .A2(_09420_),
    .ZN(_09421_));
 BUF_X4 _27784_ (.A(_09421_),
    .Z(_09422_));
 MUX2_X1 _27785_ (.A(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .B(_09419_),
    .S(_09422_),
    .Z(_02608_));
 BUF_X2 _27786_ (.A(_05409_),
    .Z(_09423_));
 MUX2_X1 _27787_ (.A(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .B(_09423_),
    .S(_09422_),
    .Z(_02609_));
 NAND2_X4 _27788_ (.A1(_04854_),
    .A2(_09420_),
    .ZN(_09424_));
 CLKBUF_X3 _27789_ (.A(_09424_),
    .Z(_09425_));
 NAND2_X1 _27790_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .A2(_09425_),
    .ZN(_09426_));
 OAI21_X1 _27791_ (.A(_09426_),
    .B1(_09425_),
    .B2(_09307_),
    .ZN(_02610_));
 NAND2_X1 _27792_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .A2(_09425_),
    .ZN(_09427_));
 OAI21_X1 _27793_ (.A(_09427_),
    .B1(_09425_),
    .B2(_09309_),
    .ZN(_02611_));
 MUX2_X1 _27794_ (.A(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .B(_09178_),
    .S(_09422_),
    .Z(_02612_));
 MUX2_X1 _27795_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .S(_09424_),
    .Z(_02613_));
 MUX2_X1 _27796_ (.A(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .B(_09180_),
    .S(_09422_),
    .Z(_02614_));
 MUX2_X1 _27797_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .S(_09424_),
    .Z(_02615_));
 NOR2_X1 _27798_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .A2(_09422_),
    .ZN(_09428_));
 AOI21_X1 _27799_ (.A(_09428_),
    .B1(_09422_),
    .B2(_09384_),
    .ZN(_02616_));
 MUX2_X1 _27800_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .S(_09424_),
    .Z(_02617_));
 NOR2_X1 _27801_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .A2(_09336_),
    .ZN(_09429_));
 AOI21_X1 _27802_ (.A(_09429_),
    .B1(_09336_),
    .B2(_09318_),
    .ZN(_02618_));
 BUF_X2 _27803_ (.A(_05761_),
    .Z(_09430_));
 BUF_X4 _27804_ (.A(_09421_),
    .Z(_09431_));
 MUX2_X1 _27805_ (.A(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .B(_09430_),
    .S(_09431_),
    .Z(_02619_));
 BUF_X2 _27806_ (.A(_05801_),
    .Z(_09432_));
 MUX2_X1 _27807_ (.A(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .B(_09432_),
    .S(_09431_),
    .Z(_02620_));
 NOR2_X1 _27808_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .A2(_09422_),
    .ZN(_09433_));
 AOI21_X1 _27809_ (.A(_09433_),
    .B1(_09422_),
    .B2(_09316_),
    .ZN(_02621_));
 MUX2_X1 _27810_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .S(_09424_),
    .Z(_02622_));
 MUX2_X1 _27811_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .S(_09424_),
    .Z(_02623_));
 BUF_X4 _27812_ (.A(_05973_),
    .Z(_09434_));
 MUX2_X1 _27813_ (.A(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .B(net403),
    .S(_09431_),
    .Z(_02624_));
 NOR2_X1 _27814_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .A2(_09422_),
    .ZN(_09435_));
 AOI21_X1 _27815_ (.A(_09435_),
    .B1(_09422_),
    .B2(_09318_),
    .ZN(_02625_));
 MUX2_X1 _27816_ (.A(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .B(_09192_),
    .S(_09431_),
    .Z(_02626_));
 MUX2_X1 _27817_ (.A(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .B(_09193_),
    .S(_09431_),
    .Z(_02627_));
 NAND2_X1 _27818_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .A2(_09425_),
    .ZN(_09436_));
 NAND2_X2 _27819_ (.A1(_05805_),
    .A2(_09420_),
    .ZN(_09437_));
 OAI21_X1 _27820_ (.A(_09436_),
    .B1(_09437_),
    .B2(_09292_),
    .ZN(_02628_));
 BUF_X2 _27821_ (.A(_06061_),
    .Z(_09438_));
 MUX2_X1 _27822_ (.A(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .B(_09438_),
    .S(_09395_),
    .Z(_02629_));
 BUF_X2 _27823_ (.A(_05543_),
    .Z(_09439_));
 MUX2_X1 _27824_ (.A(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B(_09439_),
    .S(_09236_),
    .Z(_02630_));
 MUX2_X1 _27825_ (.A(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .B(net404),
    .S(_09431_),
    .Z(_02631_));
 MUX2_X1 _27826_ (.A(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .B(_09196_),
    .S(_09431_),
    .Z(_02632_));
 MUX2_X1 _27827_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .S(_09424_),
    .Z(_02633_));
 MUX2_X1 _27828_ (.A(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .B(_09198_),
    .S(_09431_),
    .Z(_02634_));
 NAND2_X1 _27829_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A2(_09425_),
    .ZN(_09440_));
 OAI21_X1 _27830_ (.A(_09440_),
    .B1(_09437_),
    .B2(net412),
    .ZN(_02635_));
 NAND2_X1 _27831_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A2(_09425_),
    .ZN(_09441_));
 OAI21_X1 _27832_ (.A(_09441_),
    .B1(_09425_),
    .B2(_09297_),
    .ZN(_02636_));
 MUX2_X1 _27833_ (.A(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .B(net419),
    .S(_09431_),
    .Z(_02637_));
 MUX2_X1 _27834_ (.A(_09293_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .S(_09424_),
    .Z(_02638_));
 BUF_X4 _27835_ (.A(_05093_),
    .Z(_09442_));
 MUX2_X1 _27836_ (.A(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .B(net410),
    .S(_09431_),
    .Z(_02639_));
 NAND2_X1 _27837_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A2(_09425_),
    .ZN(_09443_));
 OAI21_X4 _27838_ (.A(_09443_),
    .B1(net444),
    .B2(_09437_),
    .ZN(_02640_));
 BUF_X2 _27839_ (.A(_06099_),
    .Z(_09444_));
 MUX2_X1 _27840_ (.A(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .B(_09444_),
    .S(_09395_),
    .Z(_02641_));
 BUF_X4 _27841_ (.A(_05210_),
    .Z(_09445_));
 MUX2_X1 _27842_ (.A(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .B(net356),
    .S(_09421_),
    .Z(_02642_));
 NAND2_X1 _27843_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A2(_09425_),
    .ZN(_09446_));
 OAI21_X4 _27844_ (.A(_09446_),
    .B1(net422),
    .B2(_09437_),
    .ZN(_02643_));
 AND2_X1 _27845_ (.A1(_04604_),
    .A2(_05413_),
    .ZN(_09447_));
 BUF_X4 _27846_ (.A(_09447_),
    .Z(_09448_));
 MUX2_X1 _27847_ (.A(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .B(_09419_),
    .S(_09448_),
    .Z(_02644_));
 MUX2_X1 _27848_ (.A(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .B(_09423_),
    .S(_09448_),
    .Z(_02645_));
 NAND2_X4 _27849_ (.A1(_04604_),
    .A2(_04854_),
    .ZN(_09449_));
 CLKBUF_X3 _27850_ (.A(_09449_),
    .Z(_09450_));
 NAND2_X1 _27851_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .A2(_09450_),
    .ZN(_09451_));
 OAI21_X1 _27852_ (.A(_09451_),
    .B1(_09450_),
    .B2(_09307_),
    .ZN(_02646_));
 NAND2_X1 _27853_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .A2(_09450_),
    .ZN(_09452_));
 OAI21_X1 _27854_ (.A(_09452_),
    .B1(_09450_),
    .B2(_09309_),
    .ZN(_02647_));
 MUX2_X1 _27855_ (.A(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .B(_09439_),
    .S(_09448_),
    .Z(_02648_));
 MUX2_X1 _27856_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .S(_09449_),
    .Z(_02649_));
 BUF_X2 _27857_ (.A(_05613_),
    .Z(_09453_));
 MUX2_X1 _27858_ (.A(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .B(_09453_),
    .S(_09448_),
    .Z(_02650_));
 MUX2_X1 _27859_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .S(_09449_),
    .Z(_02651_));
 NAND2_X1 _27860_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .A2(_09344_),
    .ZN(_09454_));
 NAND2_X2 _27861_ (.A1(_05805_),
    .A2(_09300_),
    .ZN(_09455_));
 OAI21_X1 _27862_ (.A(_09454_),
    .B1(_09455_),
    .B2(_09292_),
    .ZN(_02652_));
 NOR2_X1 _27863_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .A2(_09448_),
    .ZN(_09456_));
 AOI21_X1 _27864_ (.A(_09456_),
    .B1(_09448_),
    .B2(_09384_),
    .ZN(_02653_));
 MUX2_X1 _27865_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .S(_09449_),
    .Z(_02654_));
 BUF_X4 _27866_ (.A(_09447_),
    .Z(_09457_));
 MUX2_X1 _27867_ (.A(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .B(_09430_),
    .S(_09457_),
    .Z(_02655_));
 MUX2_X1 _27868_ (.A(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .B(_09432_),
    .S(_09457_),
    .Z(_02656_));
 NOR2_X1 _27869_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .A2(_09448_),
    .ZN(_09458_));
 AOI21_X1 _27870_ (.A(_09458_),
    .B1(_09448_),
    .B2(_09316_),
    .ZN(_02657_));
 MUX2_X1 _27871_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .S(_09449_),
    .Z(_02658_));
 MUX2_X1 _27872_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .S(_09449_),
    .Z(_02659_));
 MUX2_X1 _27873_ (.A(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .B(_09434_),
    .S(_09457_),
    .Z(_02660_));
 NOR2_X1 _27874_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .A2(_09448_),
    .ZN(_09459_));
 AOI21_X1 _27875_ (.A(_09459_),
    .B1(_09448_),
    .B2(_09318_),
    .ZN(_02661_));
 MUX2_X1 _27876_ (.A(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .B(_09438_),
    .S(_09457_),
    .Z(_02662_));
 BUF_X4 _27877_ (.A(_06173_),
    .Z(_09460_));
 MUX2_X1 _27878_ (.A(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .B(net406),
    .S(_09395_),
    .Z(_02663_));
 MUX2_X1 _27879_ (.A(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .B(_09444_),
    .S(_09457_),
    .Z(_02664_));
 NAND2_X1 _27880_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .A2(_09450_),
    .ZN(_09461_));
 NAND2_X2 _27881_ (.A1(_04604_),
    .A2(_05805_),
    .ZN(_09462_));
 OAI21_X1 _27882_ (.A(_09461_),
    .B1(_09462_),
    .B2(_09292_),
    .ZN(_02665_));
 MUX2_X1 _27883_ (.A(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .B(_09460_),
    .S(_09457_),
    .Z(_02666_));
 BUF_X2 _27884_ (.A(_06206_),
    .Z(_09463_));
 MUX2_X1 _27885_ (.A(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .B(_09463_),
    .S(_09457_),
    .Z(_02667_));
 MUX2_X1 _27886_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .S(_09449_),
    .Z(_02668_));
 BUF_X2 _27887_ (.A(_04765_),
    .Z(_09464_));
 MUX2_X1 _27888_ (.A(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .B(_09464_),
    .S(_09457_),
    .Z(_02669_));
 NAND2_X1 _27889_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .A2(_09450_),
    .ZN(_09465_));
 OAI21_X1 _27890_ (.A(_09465_),
    .B1(_09462_),
    .B2(net412),
    .ZN(_02670_));
 NAND2_X1 _27891_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .A2(_09450_),
    .ZN(_09466_));
 OAI21_X1 _27892_ (.A(_09466_),
    .B1(_09450_),
    .B2(_09297_),
    .ZN(_02671_));
 BUF_X4 _27893_ (.A(_05036_),
    .Z(_09467_));
 MUX2_X1 _27894_ (.A(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .B(_09467_),
    .S(_09457_),
    .Z(_02672_));
 MUX2_X1 _27895_ (.A(_09293_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .S(_09449_),
    .Z(_02673_));
 MUX2_X1 _27896_ (.A(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .B(_09463_),
    .S(_09395_),
    .Z(_02674_));
 MUX2_X1 _27897_ (.A(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .B(_09442_),
    .S(_09457_),
    .Z(_02675_));
 NAND2_X1 _27898_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .A2(_09450_),
    .ZN(_09468_));
 OAI21_X4 _27899_ (.A(_09468_),
    .B1(net444),
    .B2(_09462_),
    .ZN(_02676_));
 MUX2_X1 _27900_ (.A(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .B(_09445_),
    .S(_09447_),
    .Z(_02677_));
 NAND2_X1 _27901_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A2(_09450_),
    .ZN(_09469_));
 OAI21_X4 _27902_ (.A(_09469_),
    .B1(net422),
    .B2(_09462_),
    .ZN(_02678_));
 AND2_X1 _27903_ (.A1(_05413_),
    .A2(_05374_),
    .ZN(_09470_));
 BUF_X4 _27904_ (.A(_09470_),
    .Z(_09471_));
 MUX2_X1 _27905_ (.A(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .B(_09419_),
    .S(_09471_),
    .Z(_02679_));
 MUX2_X1 _27906_ (.A(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .B(_09423_),
    .S(_09471_),
    .Z(_02680_));
 NAND2_X4 _27907_ (.A1(_04854_),
    .A2(_05374_),
    .ZN(_09472_));
 CLKBUF_X3 _27908_ (.A(_09472_),
    .Z(_09473_));
 NAND2_X1 _27909_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .A2(_09473_),
    .ZN(_09474_));
 CLKBUF_X3 _27910_ (.A(_05463_),
    .Z(_09475_));
 OAI21_X1 _27911_ (.A(_09474_),
    .B1(_09473_),
    .B2(_09475_),
    .ZN(_02681_));
 NAND2_X1 _27912_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .A2(_09473_),
    .ZN(_09476_));
 CLKBUF_X3 _27913_ (.A(_05509_),
    .Z(_09477_));
 OAI21_X1 _27914_ (.A(_09476_),
    .B1(_09473_),
    .B2(_09477_),
    .ZN(_02682_));
 MUX2_X1 _27915_ (.A(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .B(_09439_),
    .S(_09471_),
    .Z(_02683_));
 MUX2_X1 _27916_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .S(_09472_),
    .Z(_02684_));
 MUX2_X1 _27917_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .S(_09343_),
    .Z(_02685_));
 MUX2_X1 _27918_ (.A(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .B(_09453_),
    .S(_09471_),
    .Z(_02686_));
 MUX2_X1 _27919_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .S(_09472_),
    .Z(_02687_));
 NOR2_X1 _27920_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .A2(_09471_),
    .ZN(_09478_));
 AOI21_X1 _27921_ (.A(_09478_),
    .B1(_09471_),
    .B2(_09384_),
    .ZN(_02688_));
 MUX2_X1 _27922_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .S(_09472_),
    .Z(_02689_));
 BUF_X4 _27923_ (.A(_09470_),
    .Z(_09479_));
 MUX2_X1 _27924_ (.A(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .B(_09430_),
    .S(_09479_),
    .Z(_02690_));
 MUX2_X1 _27925_ (.A(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .B(_09432_),
    .S(_09479_),
    .Z(_02691_));
 NOR2_X1 _27926_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .A2(_09471_),
    .ZN(_09480_));
 AOI21_X1 _27927_ (.A(_09480_),
    .B1(_09471_),
    .B2(_09316_),
    .ZN(_02692_));
 MUX2_X1 _27928_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .S(_09472_),
    .Z(_02693_));
 MUX2_X1 _27929_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .S(_09472_),
    .Z(_02694_));
 MUX2_X1 _27930_ (.A(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .B(net403),
    .S(_09479_),
    .Z(_02695_));
 MUX2_X1 _27931_ (.A(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .B(_09464_),
    .S(_09395_),
    .Z(_02696_));
 NOR2_X1 _27932_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .A2(_09471_),
    .ZN(_09481_));
 AOI21_X1 _27933_ (.A(_09481_),
    .B1(_09471_),
    .B2(_09318_),
    .ZN(_02697_));
 MUX2_X1 _27934_ (.A(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .B(_09438_),
    .S(_09479_),
    .Z(_02698_));
 MUX2_X1 _27935_ (.A(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .B(_09444_),
    .S(_09479_),
    .Z(_02699_));
 NAND2_X1 _27936_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .A2(_09473_),
    .ZN(_09482_));
 NAND2_X2 _27937_ (.A1(_05805_),
    .A2(_05374_),
    .ZN(_09483_));
 CLKBUF_X3 _27938_ (.A(_06137_),
    .Z(_09484_));
 OAI21_X1 _27939_ (.A(_09482_),
    .B1(_09483_),
    .B2(_09484_),
    .ZN(_02700_));
 MUX2_X1 _27940_ (.A(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .B(net406),
    .S(_09479_),
    .Z(_02701_));
 MUX2_X1 _27941_ (.A(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .B(_09463_),
    .S(_09479_),
    .Z(_02702_));
 MUX2_X1 _27942_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .S(_09472_),
    .Z(_02703_));
 MUX2_X1 _27943_ (.A(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .B(_09464_),
    .S(_09479_),
    .Z(_02704_));
 NAND2_X1 _27944_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .A2(_09473_),
    .ZN(_09485_));
 OAI21_X1 _27945_ (.A(_09485_),
    .B1(_09483_),
    .B2(net412),
    .ZN(_02705_));
 NAND2_X1 _27946_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .A2(_09473_),
    .ZN(_09486_));
 OAI21_X1 _27947_ (.A(_09486_),
    .B1(_09473_),
    .B2(_09297_),
    .ZN(_02706_));
 NAND2_X1 _27948_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A2(_09344_),
    .ZN(_09487_));
 BUF_X8 _27949_ (.A(_04907_),
    .Z(_09488_));
 OAI21_X1 _27950_ (.A(_09487_),
    .B1(_09455_),
    .B2(_09488_),
    .ZN(_02707_));
 MUX2_X1 _27951_ (.A(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .B(_09467_),
    .S(_09479_),
    .Z(_02708_));
 MUX2_X1 _27952_ (.A(_09293_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .S(_09472_),
    .Z(_02709_));
 MUX2_X1 _27953_ (.A(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .B(_09442_),
    .S(_09479_),
    .Z(_02710_));
 NAND2_X1 _27954_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .A2(_09473_),
    .ZN(_09489_));
 OAI21_X4 _27955_ (.A(_09489_),
    .B1(net444),
    .B2(_09483_),
    .ZN(_02711_));
 MUX2_X1 _27956_ (.A(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .B(net356),
    .S(_09470_),
    .Z(_02712_));
 NAND2_X1 _27957_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A2(_09473_),
    .ZN(_09490_));
 OAI21_X4 _27958_ (.A(_09490_),
    .B1(net422),
    .B2(_09483_),
    .ZN(_02713_));
 AND2_X1 _27959_ (.A1(_05413_),
    .A2(_06214_),
    .ZN(_09491_));
 BUF_X4 _27960_ (.A(_09491_),
    .Z(_09492_));
 MUX2_X1 _27961_ (.A(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .B(_09419_),
    .S(_09492_),
    .Z(_02714_));
 MUX2_X1 _27962_ (.A(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .B(_09423_),
    .S(_09492_),
    .Z(_02715_));
 NAND2_X4 _27963_ (.A1(_04854_),
    .A2(_06214_),
    .ZN(_09493_));
 CLKBUF_X3 _27964_ (.A(_09493_),
    .Z(_09494_));
 NAND2_X1 _27965_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .A2(_09494_),
    .ZN(_09495_));
 OAI21_X1 _27966_ (.A(_09495_),
    .B1(_09494_),
    .B2(_09475_),
    .ZN(_02716_));
 NAND2_X1 _27967_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .A2(_09494_),
    .ZN(_09496_));
 OAI21_X1 _27968_ (.A(_09496_),
    .B1(_09494_),
    .B2(_09477_),
    .ZN(_02717_));
 NAND2_X1 _27969_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .A2(_09344_),
    .ZN(_09497_));
 BUF_X8 _27970_ (.A(_04977_),
    .Z(_09498_));
 OAI21_X1 _27971_ (.A(_09497_),
    .B1(_09344_),
    .B2(_09498_),
    .ZN(_02718_));
 MUX2_X1 _27972_ (.A(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .B(_09439_),
    .S(_09492_),
    .Z(_02719_));
 MUX2_X1 _27973_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S(_09493_),
    .Z(_02720_));
 MUX2_X1 _27974_ (.A(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .B(_09453_),
    .S(_09492_),
    .Z(_02721_));
 MUX2_X1 _27975_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(_09493_),
    .Z(_02722_));
 NOR2_X1 _27976_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .A2(_09492_),
    .ZN(_09499_));
 AOI21_X1 _27977_ (.A(_09499_),
    .B1(_09492_),
    .B2(_09384_),
    .ZN(_02723_));
 MUX2_X1 _27978_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S(_09493_),
    .Z(_02724_));
 BUF_X4 _27979_ (.A(_09491_),
    .Z(_09500_));
 MUX2_X1 _27980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .B(_09430_),
    .S(_09500_),
    .Z(_02725_));
 MUX2_X1 _27981_ (.A(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .B(_09432_),
    .S(_09500_),
    .Z(_02726_));
 NOR2_X1 _27982_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .A2(_09492_),
    .ZN(_09501_));
 AOI21_X1 _27983_ (.A(_09501_),
    .B1(_09492_),
    .B2(_09316_),
    .ZN(_02727_));
 MUX2_X1 _27984_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(_09493_),
    .Z(_02728_));
 MUX2_X1 _27985_ (.A(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .B(_09467_),
    .S(_09395_),
    .Z(_02729_));
 MUX2_X1 _27986_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(_09493_),
    .Z(_02730_));
 MUX2_X1 _27987_ (.A(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .B(net403),
    .S(_09500_),
    .Z(_02731_));
 NOR2_X1 _27988_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .A2(_09492_),
    .ZN(_09502_));
 AOI21_X1 _27989_ (.A(_09502_),
    .B1(_09492_),
    .B2(_09318_),
    .ZN(_02732_));
 MUX2_X1 _27990_ (.A(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .B(_09438_),
    .S(_09500_),
    .Z(_02733_));
 MUX2_X1 _27991_ (.A(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .B(_09444_),
    .S(_09500_),
    .Z(_02734_));
 NAND2_X1 _27992_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .A2(_09494_),
    .ZN(_09503_));
 NAND2_X2 _27993_ (.A1(_05805_),
    .A2(_06214_),
    .ZN(_09504_));
 OAI21_X1 _27994_ (.A(_09503_),
    .B1(_09504_),
    .B2(_09484_),
    .ZN(_02735_));
 MUX2_X1 _27995_ (.A(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .B(_09460_),
    .S(_09500_),
    .Z(_02736_));
 MUX2_X1 _27996_ (.A(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .B(_09463_),
    .S(_09500_),
    .Z(_02737_));
 MUX2_X1 _27997_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S(_09493_),
    .Z(_02738_));
 MUX2_X1 _27998_ (.A(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .B(_09464_),
    .S(_09500_),
    .Z(_02739_));
 MUX2_X1 _27999_ (.A(net332),
    .B(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .S(_09343_),
    .Z(_02740_));
 MUX2_X1 _28000_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .S(_06246_),
    .Z(_02741_));
 NAND2_X1 _28001_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .A2(_09494_),
    .ZN(_09505_));
 OAI21_X1 _28002_ (.A(_09505_),
    .B1(_09504_),
    .B2(net420),
    .ZN(_02742_));
 NAND2_X1 _28003_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .A2(_09494_),
    .ZN(_09506_));
 OAI21_X1 _28004_ (.A(_09506_),
    .B1(_09494_),
    .B2(_09498_),
    .ZN(_02743_));
 MUX2_X1 _28005_ (.A(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .B(net440),
    .S(_09500_),
    .Z(_02744_));
 MUX2_X1 _28006_ (.A(net332),
    .B(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S(_09493_),
    .Z(_02745_));
 MUX2_X1 _28007_ (.A(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .B(_09442_),
    .S(_09500_),
    .Z(_02746_));
 NAND2_X1 _28008_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .A2(_09494_),
    .ZN(_09507_));
 BUF_X16 _28009_ (.A(_05147_),
    .Z(_09508_));
 OAI21_X4 _28010_ (.A(_09507_),
    .B1(net447),
    .B2(_09504_),
    .ZN(_02747_));
 MUX2_X1 _28011_ (.A(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .B(_09445_),
    .S(_09491_),
    .Z(_02748_));
 NAND2_X1 _28012_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .A2(_09494_),
    .ZN(_09509_));
 BUF_X8 _28013_ (.A(_05259_),
    .Z(_09510_));
 OAI21_X4 _28014_ (.A(_09509_),
    .B1(net438),
    .B2(_09504_),
    .ZN(_02749_));
 AND3_X1 _28015_ (.A1(_05412_),
    .A2(_06226_),
    .A3(_09420_),
    .ZN(_09511_));
 BUF_X4 _28016_ (.A(_09511_),
    .Z(_09512_));
 BUF_X4 _28017_ (.A(_09512_),
    .Z(_09513_));
 MUX2_X1 _28018_ (.A(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .B(_09419_),
    .S(_09513_),
    .Z(_02750_));
 MUX2_X1 _28019_ (.A(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .B(_09423_),
    .S(_09513_),
    .Z(_02751_));
 MUX2_X1 _28020_ (.A(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .B(net410),
    .S(_09395_),
    .Z(_02752_));
 NAND3_X4 _28021_ (.A1(_06224_),
    .A2(_06226_),
    .A3(_09420_),
    .ZN(_09514_));
 CLKBUF_X3 _28022_ (.A(_09514_),
    .Z(_09515_));
 NAND2_X1 _28023_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .A2(_09515_),
    .ZN(_09516_));
 OAI21_X1 _28024_ (.A(_09516_),
    .B1(_09515_),
    .B2(_09475_),
    .ZN(_02753_));
 NAND2_X1 _28025_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .A2(_09515_),
    .ZN(_09517_));
 OAI21_X1 _28026_ (.A(_09517_),
    .B1(_09515_),
    .B2(_09477_),
    .ZN(_02754_));
 MUX2_X1 _28027_ (.A(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .B(_09439_),
    .S(_09513_),
    .Z(_02755_));
 MUX2_X1 _28028_ (.A(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .B(_09179_),
    .S(_09513_),
    .Z(_02756_));
 MUX2_X1 _28029_ (.A(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .B(_09453_),
    .S(_09513_),
    .Z(_02757_));
 MUX2_X1 _28030_ (.A(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .B(_09181_),
    .S(_09513_),
    .Z(_02758_));
 NAND2_X1 _28031_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .A2(_09514_),
    .ZN(_09518_));
 OAI21_X1 _28032_ (.A(_09518_),
    .B1(_09515_),
    .B2(_06222_),
    .ZN(_02759_));
 BUF_X4 _28033_ (.A(_09512_),
    .Z(_09519_));
 MUX2_X1 _28034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .B(_09183_),
    .S(_09519_),
    .Z(_02760_));
 MUX2_X1 _28035_ (.A(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .B(_09430_),
    .S(_09519_),
    .Z(_02761_));
 MUX2_X1 _28036_ (.A(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .B(_09432_),
    .S(_09519_),
    .Z(_02762_));
 NAND2_X1 _28037_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A2(_09344_),
    .ZN(_09520_));
 OAI21_X1 _28038_ (.A(_09520_),
    .B1(_09455_),
    .B2(_09508_),
    .ZN(_02763_));
 NOR2_X1 _28039_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .A2(_09513_),
    .ZN(_09521_));
 AOI21_X1 _28040_ (.A(_09521_),
    .B1(_09513_),
    .B2(_09316_),
    .ZN(_02764_));
 MUX2_X1 _28041_ (.A(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .B(_09188_),
    .S(_09519_),
    .Z(_02765_));
 MUX2_X1 _28042_ (.A(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .B(_09189_),
    .S(_09519_),
    .Z(_02766_));
 MUX2_X1 _28043_ (.A(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .B(_09434_),
    .S(_09519_),
    .Z(_02767_));
 NOR2_X1 _28044_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .A2(_09513_),
    .ZN(_09522_));
 AOI21_X1 _28045_ (.A(_09522_),
    .B1(_09513_),
    .B2(_09318_),
    .ZN(_02768_));
 MUX2_X1 _28046_ (.A(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .B(_09438_),
    .S(_09519_),
    .Z(_02769_));
 MUX2_X1 _28047_ (.A(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .B(_09444_),
    .S(_09519_),
    .Z(_02770_));
 NAND2_X1 _28048_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .A2(_09514_),
    .ZN(_09523_));
 OAI21_X1 _28049_ (.A(_09523_),
    .B1(_09515_),
    .B2(_09484_),
    .ZN(_02771_));
 MUX2_X1 _28050_ (.A(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .B(_09460_),
    .S(_09519_),
    .Z(_02772_));
 MUX2_X1 _28051_ (.A(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .B(_09463_),
    .S(_09519_),
    .Z(_02773_));
 MUX2_X1 _28052_ (.A(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .B(_09445_),
    .S(_09335_),
    .Z(_02774_));
 MUX2_X1 _28053_ (.A(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .B(_09197_),
    .S(_09512_),
    .Z(_02775_));
 MUX2_X1 _28054_ (.A(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .B(_09464_),
    .S(_09512_),
    .Z(_02776_));
 NAND2_X1 _28055_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A2(_09514_),
    .ZN(_09524_));
 OAI21_X1 _28056_ (.A(_09524_),
    .B1(_09515_),
    .B2(_09488_),
    .ZN(_02777_));
 NAND2_X1 _28057_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A2(_09514_),
    .ZN(_09525_));
 OAI21_X1 _28058_ (.A(_09525_),
    .B1(_09515_),
    .B2(_09498_),
    .ZN(_02778_));
 MUX2_X1 _28059_ (.A(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .B(_09467_),
    .S(_09512_),
    .Z(_02779_));
 MUX2_X1 _28060_ (.A(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .B(_09202_),
    .S(_09512_),
    .Z(_02780_));
 MUX2_X1 _28061_ (.A(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .B(_09442_),
    .S(_09512_),
    .Z(_02781_));
 NAND2_X1 _28062_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A2(_09514_),
    .ZN(_09526_));
 OAI21_X4 _28063_ (.A(_09526_),
    .B1(net447),
    .B2(_09515_),
    .ZN(_02782_));
 MUX2_X1 _28064_ (.A(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .B(net356),
    .S(_09512_),
    .Z(_02783_));
 NAND2_X1 _28065_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A2(_09514_),
    .ZN(_09527_));
 OAI21_X4 _28066_ (.A(_09527_),
    .B1(net438),
    .B2(_09515_),
    .ZN(_02784_));
 NAND2_X1 _28067_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(_09344_),
    .ZN(_09528_));
 OAI21_X4 _28068_ (.A(_09528_),
    .B1(net438),
    .B2(_09455_),
    .ZN(_02785_));
 AND3_X1 _28069_ (.A1(_05412_),
    .A2(_04604_),
    .A3(_06225_),
    .ZN(_09529_));
 BUF_X4 _28070_ (.A(_09529_),
    .Z(_09530_));
 BUF_X4 _28071_ (.A(_09530_),
    .Z(_09531_));
 MUX2_X1 _28072_ (.A(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .B(_09419_),
    .S(_09531_),
    .Z(_02786_));
 MUX2_X1 _28073_ (.A(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .B(_09423_),
    .S(_09531_),
    .Z(_02787_));
 NAND3_X2 _28074_ (.A1(_06224_),
    .A2(_04604_),
    .A3(_06226_),
    .ZN(_09532_));
 CLKBUF_X3 _28075_ (.A(_09532_),
    .Z(_09533_));
 NAND2_X1 _28076_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .A2(_09533_),
    .ZN(_09534_));
 OAI21_X1 _28077_ (.A(_09534_),
    .B1(_09533_),
    .B2(_09475_),
    .ZN(_02788_));
 NAND2_X1 _28078_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .A2(_09533_),
    .ZN(_09535_));
 OAI21_X1 _28079_ (.A(_09535_),
    .B1(_09533_),
    .B2(_09477_),
    .ZN(_02789_));
 MUX2_X1 _28080_ (.A(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .B(_09439_),
    .S(_09531_),
    .Z(_02790_));
 MUX2_X1 _28081_ (.A(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .B(_09179_),
    .S(_09531_),
    .Z(_02791_));
 BUF_X4 _28082_ (.A(_09530_),
    .Z(_09536_));
 MUX2_X1 _28083_ (.A(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .B(_09453_),
    .S(_09536_),
    .Z(_02792_));
 MUX2_X1 _28084_ (.A(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .B(_09181_),
    .S(_09536_),
    .Z(_02793_));
 NOR2_X1 _28085_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .A2(_09531_),
    .ZN(_09537_));
 AOI21_X1 _28086_ (.A(_09537_),
    .B1(_09531_),
    .B2(_09384_),
    .ZN(_02794_));
 MUX2_X1 _28087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .B(_09183_),
    .S(_09536_),
    .Z(_02795_));
 MUX2_X1 _28088_ (.A(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .B(_09419_),
    .S(_05415_),
    .Z(_02796_));
 MUX2_X1 _28089_ (.A(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .B(_09430_),
    .S(_09536_),
    .Z(_02797_));
 MUX2_X1 _28090_ (.A(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .B(_09432_),
    .S(_09536_),
    .Z(_02798_));
 NOR2_X1 _28091_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .A2(_09531_),
    .ZN(_09538_));
 AOI21_X1 _28092_ (.A(_09538_),
    .B1(_09531_),
    .B2(_09316_),
    .ZN(_02799_));
 MUX2_X1 _28093_ (.A(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .B(_09188_),
    .S(_09536_),
    .Z(_02800_));
 MUX2_X1 _28094_ (.A(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .B(_09189_),
    .S(_09536_),
    .Z(_02801_));
 MUX2_X1 _28095_ (.A(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .B(_09434_),
    .S(_09536_),
    .Z(_02802_));
 NOR2_X1 _28096_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .A2(_09531_),
    .ZN(_09539_));
 AOI21_X1 _28097_ (.A(_09539_),
    .B1(_09531_),
    .B2(_09318_),
    .ZN(_02803_));
 MUX2_X1 _28098_ (.A(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .B(_09438_),
    .S(_09536_),
    .Z(_02804_));
 MUX2_X1 _28099_ (.A(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .B(_09444_),
    .S(_09536_),
    .Z(_02805_));
 NAND2_X1 _28100_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .A2(_09533_),
    .ZN(_09540_));
 OAI21_X1 _28101_ (.A(_09540_),
    .B1(_09533_),
    .B2(_09484_),
    .ZN(_02806_));
 MUX2_X1 _28102_ (.A(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .B(_09423_),
    .S(_05415_),
    .Z(_02807_));
 MUX2_X1 _28103_ (.A(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .B(net406),
    .S(_09530_),
    .Z(_02808_));
 MUX2_X1 _28104_ (.A(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .B(_09463_),
    .S(_09530_),
    .Z(_02809_));
 MUX2_X1 _28105_ (.A(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .B(_09197_),
    .S(_09530_),
    .Z(_02810_));
 MUX2_X1 _28106_ (.A(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .B(_09464_),
    .S(_09530_),
    .Z(_02811_));
 NAND2_X1 _28107_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .A2(_09532_),
    .ZN(_09541_));
 OAI21_X1 _28108_ (.A(_09541_),
    .B1(_09533_),
    .B2(net420),
    .ZN(_02812_));
 NAND2_X1 _28109_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .A2(_09532_),
    .ZN(_09542_));
 OAI21_X1 _28110_ (.A(_09542_),
    .B1(_09533_),
    .B2(_09498_),
    .ZN(_02813_));
 MUX2_X1 _28111_ (.A(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .B(net440),
    .S(_09530_),
    .Z(_02814_));
 MUX2_X1 _28112_ (.A(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .B(_09202_),
    .S(_09530_),
    .Z(_02815_));
 MUX2_X1 _28113_ (.A(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .B(net410),
    .S(_09530_),
    .Z(_02816_));
 NAND2_X1 _28114_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .A2(_09532_),
    .ZN(_09543_));
 OAI21_X4 _28115_ (.A(_09543_),
    .B1(net447),
    .B2(_09533_),
    .ZN(_02817_));
 NAND2_X1 _28116_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .A2(_05803_),
    .ZN(_09544_));
 OAI21_X1 _28117_ (.A(_09544_),
    .B1(_05464_),
    .B2(_05803_),
    .ZN(_02818_));
 MUX2_X1 _28118_ (.A(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .B(net356),
    .S(_09530_),
    .Z(_02819_));
 NAND2_X1 _28119_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A2(_09532_),
    .ZN(_09545_));
 OAI21_X4 _28120_ (.A(_09545_),
    .B1(net438),
    .B2(_09533_),
    .ZN(_02820_));
 AND3_X1 _28121_ (.A1(_05412_),
    .A2(_06225_),
    .A3(_05374_),
    .ZN(_09546_));
 BUF_X4 _28122_ (.A(_09546_),
    .Z(_09547_));
 BUF_X4 _28123_ (.A(_09547_),
    .Z(_09548_));
 MUX2_X1 _28124_ (.A(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .B(_09419_),
    .S(_09548_),
    .Z(_02821_));
 MUX2_X1 _28125_ (.A(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .B(_09423_),
    .S(_09548_),
    .Z(_02822_));
 NAND3_X2 _28126_ (.A1(_06224_),
    .A2(_06226_),
    .A3(_05374_),
    .ZN(_09549_));
 CLKBUF_X3 _28127_ (.A(_09549_),
    .Z(_09550_));
 NAND2_X1 _28128_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .A2(_09550_),
    .ZN(_09551_));
 OAI21_X1 _28129_ (.A(_09551_),
    .B1(_09550_),
    .B2(_09475_),
    .ZN(_02823_));
 NAND2_X1 _28130_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .A2(_09550_),
    .ZN(_09552_));
 OAI21_X1 _28131_ (.A(_09552_),
    .B1(_09550_),
    .B2(_09477_),
    .ZN(_02824_));
 MUX2_X1 _28132_ (.A(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .B(_09439_),
    .S(_09548_),
    .Z(_02825_));
 MUX2_X1 _28133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .B(_05580_),
    .S(_09548_),
    .Z(_02826_));
 BUF_X4 _28134_ (.A(_09547_),
    .Z(_09553_));
 MUX2_X1 _28135_ (.A(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .B(_09453_),
    .S(_09553_),
    .Z(_02827_));
 MUX2_X1 _28136_ (.A(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .B(_05653_),
    .S(_09553_),
    .Z(_02828_));
 NAND2_X1 _28137_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .A2(_05803_),
    .ZN(_09554_));
 OAI21_X1 _28138_ (.A(_09554_),
    .B1(_05510_),
    .B2(_05803_),
    .ZN(_02829_));
 NOR2_X1 _28139_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .A2(_09548_),
    .ZN(_09555_));
 AOI21_X1 _28140_ (.A(_09555_),
    .B1(_09548_),
    .B2(_09384_),
    .ZN(_02830_));
 MUX2_X1 _28141_ (.A(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .B(_05721_),
    .S(_09553_),
    .Z(_02831_));
 MUX2_X1 _28142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .B(_09430_),
    .S(_09553_),
    .Z(_02832_));
 MUX2_X1 _28143_ (.A(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .B(_09432_),
    .S(_09553_),
    .Z(_02833_));
 NOR2_X1 _28144_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .A2(_09548_),
    .ZN(_09556_));
 AOI21_X1 _28145_ (.A(_09556_),
    .B1(_09548_),
    .B2(_09316_),
    .ZN(_02834_));
 MUX2_X1 _28146_ (.A(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .B(_05890_),
    .S(_09553_),
    .Z(_02835_));
 MUX2_X1 _28147_ (.A(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .B(_05928_),
    .S(_09553_),
    .Z(_02836_));
 MUX2_X1 _28148_ (.A(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .B(net403),
    .S(_09553_),
    .Z(_02837_));
 NOR2_X1 _28149_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .A2(_09548_),
    .ZN(_09557_));
 AOI21_X1 _28150_ (.A(_09557_),
    .B1(_09548_),
    .B2(_09318_),
    .ZN(_02838_));
 MUX2_X1 _28151_ (.A(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .B(_09438_),
    .S(_09553_),
    .Z(_02839_));
 BUF_X4 _28152_ (.A(_05414_),
    .Z(_09558_));
 MUX2_X1 _28153_ (.A(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .B(_09439_),
    .S(_09558_),
    .Z(_02840_));
 MUX2_X1 _28154_ (.A(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .B(_09444_),
    .S(_09553_),
    .Z(_02841_));
 NAND2_X1 _28155_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .A2(_09550_),
    .ZN(_09559_));
 OAI21_X1 _28156_ (.A(_09559_),
    .B1(_09550_),
    .B2(_09484_),
    .ZN(_02842_));
 MUX2_X1 _28157_ (.A(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .B(net406),
    .S(_09547_),
    .Z(_02843_));
 MUX2_X1 _28158_ (.A(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .B(_09463_),
    .S(_09547_),
    .Z(_02844_));
 MUX2_X1 _28159_ (.A(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .B(_04602_),
    .S(_09547_),
    .Z(_02845_));
 MUX2_X1 _28160_ (.A(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .B(_09464_),
    .S(_09547_),
    .Z(_02846_));
 NAND2_X1 _28161_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .A2(_09549_),
    .ZN(_09560_));
 OAI21_X1 _28162_ (.A(_09560_),
    .B1(_09550_),
    .B2(_09488_),
    .ZN(_02847_));
 NAND2_X1 _28163_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .A2(_09549_),
    .ZN(_09561_));
 OAI21_X1 _28164_ (.A(_09561_),
    .B1(_09550_),
    .B2(_09498_),
    .ZN(_02848_));
 MUX2_X1 _28165_ (.A(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .B(net440),
    .S(_09547_),
    .Z(_02849_));
 MUX2_X1 _28166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .B(_04850_),
    .S(_09547_),
    .Z(_02850_));
 MUX2_X1 _28167_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(_04855_),
    .Z(_02851_));
 MUX2_X1 _28168_ (.A(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .B(_09453_),
    .S(_09176_),
    .Z(_02852_));
 MUX2_X1 _28169_ (.A(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .B(_09442_),
    .S(_09547_),
    .Z(_02853_));
 NAND2_X1 _28170_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .A2(_09549_),
    .ZN(_09562_));
 OAI21_X4 _28171_ (.A(_09562_),
    .B1(net447),
    .B2(_09550_),
    .ZN(_02854_));
 MUX2_X1 _28172_ (.A(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .B(_09445_),
    .S(_09547_),
    .Z(_02855_));
 NAND2_X1 _28173_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A2(_09549_),
    .ZN(_09563_));
 OAI21_X4 _28174_ (.A(_09563_),
    .B1(_09510_),
    .B2(_09550_),
    .ZN(_02856_));
 AND3_X1 _28175_ (.A1(_05412_),
    .A2(_06225_),
    .A3(_06214_),
    .ZN(_09564_));
 BUF_X4 _28176_ (.A(_09564_),
    .Z(_09565_));
 BUF_X4 _28177_ (.A(_09565_),
    .Z(_09566_));
 MUX2_X1 _28178_ (.A(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .B(_09419_),
    .S(_09566_),
    .Z(_02857_));
 MUX2_X1 _28179_ (.A(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .B(_09423_),
    .S(_09566_),
    .Z(_02858_));
 NAND3_X2 _28180_ (.A1(_06224_),
    .A2(_06226_),
    .A3(_06214_),
    .ZN(_09567_));
 CLKBUF_X3 _28181_ (.A(_09567_),
    .Z(_09568_));
 NAND2_X1 _28182_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .A2(_09568_),
    .ZN(_09569_));
 OAI21_X1 _28183_ (.A(_09569_),
    .B1(_09568_),
    .B2(_09475_),
    .ZN(_02859_));
 NAND2_X1 _28184_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .A2(_09568_),
    .ZN(_09570_));
 OAI21_X1 _28185_ (.A(_09570_),
    .B1(_09568_),
    .B2(_09477_),
    .ZN(_02860_));
 MUX2_X1 _28186_ (.A(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .B(_09439_),
    .S(_09566_),
    .Z(_02861_));
 MUX2_X1 _28187_ (.A(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .B(_05580_),
    .S(_09566_),
    .Z(_02862_));
 MUX2_X1 _28188_ (.A(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .B(_09453_),
    .S(_09558_),
    .Z(_02863_));
 BUF_X4 _28189_ (.A(_09565_),
    .Z(_09571_));
 MUX2_X1 _28190_ (.A(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .B(_09453_),
    .S(_09571_),
    .Z(_02864_));
 MUX2_X1 _28191_ (.A(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .B(_05653_),
    .S(_09571_),
    .Z(_02865_));
 NOR2_X1 _28192_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .A2(_09566_),
    .ZN(_09572_));
 AOI21_X1 _28193_ (.A(_09572_),
    .B1(_09566_),
    .B2(_09384_),
    .ZN(_02866_));
 MUX2_X1 _28194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .B(_05721_),
    .S(_09571_),
    .Z(_02867_));
 MUX2_X1 _28195_ (.A(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .B(_09430_),
    .S(_09571_),
    .Z(_02868_));
 MUX2_X1 _28196_ (.A(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .B(_09432_),
    .S(_09571_),
    .Z(_02869_));
 NOR2_X1 _28197_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .A2(_09566_),
    .ZN(_09573_));
 AOI21_X1 _28198_ (.A(_09573_),
    .B1(_09566_),
    .B2(_06231_),
    .ZN(_02870_));
 MUX2_X1 _28199_ (.A(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .B(_05890_),
    .S(_09571_),
    .Z(_02871_));
 MUX2_X1 _28200_ (.A(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .B(_05928_),
    .S(_09571_),
    .Z(_02872_));
 MUX2_X1 _28201_ (.A(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .B(net403),
    .S(_09571_),
    .Z(_02873_));
 MUX2_X1 _28202_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(_04855_),
    .Z(_02874_));
 NOR2_X1 _28203_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .A2(_09566_),
    .ZN(_09574_));
 AOI21_X1 _28204_ (.A(_09574_),
    .B1(_09566_),
    .B2(_06234_),
    .ZN(_02875_));
 MUX2_X1 _28205_ (.A(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .B(_09438_),
    .S(_09571_),
    .Z(_02876_));
 MUX2_X1 _28206_ (.A(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .B(_09444_),
    .S(_09571_),
    .Z(_02877_));
 NAND2_X1 _28207_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .A2(_09568_),
    .ZN(_09575_));
 OAI21_X1 _28208_ (.A(_09575_),
    .B1(_09568_),
    .B2(_09484_),
    .ZN(_02878_));
 MUX2_X1 _28209_ (.A(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .B(net406),
    .S(_09565_),
    .Z(_02879_));
 MUX2_X1 _28210_ (.A(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .B(_09463_),
    .S(_09565_),
    .Z(_02880_));
 MUX2_X1 _28211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .B(_04602_),
    .S(_09565_),
    .Z(_02881_));
 MUX2_X1 _28212_ (.A(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .B(_09464_),
    .S(_09565_),
    .Z(_02882_));
 NAND2_X1 _28213_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .A2(_09567_),
    .ZN(_09576_));
 OAI21_X1 _28214_ (.A(_09576_),
    .B1(_09568_),
    .B2(_09488_),
    .ZN(_02883_));
 NAND2_X1 _28215_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .A2(_09567_),
    .ZN(_09577_));
 OAI21_X1 _28216_ (.A(_09577_),
    .B1(_09568_),
    .B2(_09498_),
    .ZN(_02884_));
 NOR2_X1 _28217_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .A2(_05415_),
    .ZN(_09578_));
 AOI21_X1 _28218_ (.A(_09578_),
    .B1(_05688_),
    .B2(_05415_),
    .ZN(_02885_));
 MUX2_X1 _28219_ (.A(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .B(net440),
    .S(_09565_),
    .Z(_02886_));
 MUX2_X1 _28220_ (.A(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .B(_04850_),
    .S(_09565_),
    .Z(_02887_));
 MUX2_X1 _28221_ (.A(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .B(net410),
    .S(_09565_),
    .Z(_02888_));
 NAND2_X1 _28222_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .A2(_09567_),
    .ZN(_09579_));
 OAI21_X4 _28223_ (.A(_09579_),
    .B1(_09508_),
    .B2(_09568_),
    .ZN(_02889_));
 MUX2_X1 _28224_ (.A(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .B(net356),
    .S(_09565_),
    .Z(_02890_));
 NAND2_X1 _28225_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .A2(_09567_),
    .ZN(_09580_));
 OAI21_X4 _28226_ (.A(_09580_),
    .B1(_09510_),
    .B2(_09568_),
    .ZN(_02891_));
 AND2_X1 _28227_ (.A1(_09264_),
    .A2(_09420_),
    .ZN(_09581_));
 BUF_X4 _28228_ (.A(_09581_),
    .Z(_09582_));
 BUF_X4 _28229_ (.A(_09582_),
    .Z(_09583_));
 MUX2_X1 _28230_ (.A(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .B(_09419_),
    .S(_09583_),
    .Z(_02892_));
 MUX2_X1 _28231_ (.A(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .B(_09423_),
    .S(_09583_),
    .Z(_02893_));
 NAND2_X2 _28232_ (.A1(_09264_),
    .A2(_09420_),
    .ZN(_09584_));
 CLKBUF_X3 _28233_ (.A(_09584_),
    .Z(_09585_));
 NAND2_X1 _28234_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .A2(_09585_),
    .ZN(_09586_));
 OAI21_X1 _28235_ (.A(_09586_),
    .B1(_09585_),
    .B2(_09475_),
    .ZN(_02894_));
 NAND2_X1 _28236_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .A2(_09585_),
    .ZN(_09587_));
 OAI21_X1 _28237_ (.A(_09587_),
    .B1(_09585_),
    .B2(_09477_),
    .ZN(_02895_));
 MUX2_X1 _28238_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(_04855_),
    .Z(_02896_));
 MUX2_X1 _28239_ (.A(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .B(_09439_),
    .S(_09583_),
    .Z(_02897_));
 MUX2_X1 _28240_ (.A(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .B(_05580_),
    .S(_09583_),
    .Z(_02898_));
 BUF_X4 _28241_ (.A(_09582_),
    .Z(_09588_));
 MUX2_X1 _28242_ (.A(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .B(_09453_),
    .S(_09588_),
    .Z(_02899_));
 MUX2_X1 _28243_ (.A(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .B(_05653_),
    .S(_09588_),
    .Z(_02900_));
 NOR2_X1 _28244_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .A2(_09583_),
    .ZN(_09589_));
 AOI21_X1 _28245_ (.A(_09589_),
    .B1(_09583_),
    .B2(_09384_),
    .ZN(_02901_));
 MUX2_X1 _28246_ (.A(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .B(_05721_),
    .S(_09588_),
    .Z(_02902_));
 MUX2_X1 _28247_ (.A(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .B(_09430_),
    .S(_09588_),
    .Z(_02903_));
 MUX2_X1 _28248_ (.A(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .B(_09432_),
    .S(_09588_),
    .Z(_02904_));
 NOR2_X1 _28249_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .A2(_09583_),
    .ZN(_09590_));
 AOI21_X1 _28250_ (.A(_09590_),
    .B1(_09583_),
    .B2(_06231_),
    .ZN(_02905_));
 MUX2_X1 _28251_ (.A(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .B(_05890_),
    .S(_09588_),
    .Z(_02906_));
 MUX2_X1 _28252_ (.A(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .B(_09430_),
    .S(_09558_),
    .Z(_02907_));
 MUX2_X1 _28253_ (.A(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .B(_05928_),
    .S(_09588_),
    .Z(_02908_));
 MUX2_X1 _28254_ (.A(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .B(_09434_),
    .S(_09588_),
    .Z(_02909_));
 NOR2_X1 _28255_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .A2(_09583_),
    .ZN(_09591_));
 AOI21_X1 _28256_ (.A(_09591_),
    .B1(_09583_),
    .B2(_06234_),
    .ZN(_02910_));
 MUX2_X1 _28257_ (.A(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .B(_09438_),
    .S(_09588_),
    .Z(_02911_));
 MUX2_X1 _28258_ (.A(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .B(_09444_),
    .S(_09588_),
    .Z(_02912_));
 NAND2_X1 _28259_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .A2(_09585_),
    .ZN(_09592_));
 OAI21_X1 _28260_ (.A(_09592_),
    .B1(_09585_),
    .B2(_09484_),
    .ZN(_02913_));
 MUX2_X1 _28261_ (.A(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .B(_09460_),
    .S(_09582_),
    .Z(_02914_));
 MUX2_X1 _28262_ (.A(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .B(_09463_),
    .S(_09582_),
    .Z(_02915_));
 MUX2_X1 _28263_ (.A(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .B(_04602_),
    .S(_09582_),
    .Z(_02916_));
 MUX2_X1 _28264_ (.A(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .B(_09464_),
    .S(_09582_),
    .Z(_02917_));
 MUX2_X1 _28265_ (.A(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .B(_09432_),
    .S(_09558_),
    .Z(_02918_));
 NAND2_X1 _28266_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A2(_09584_),
    .ZN(_09593_));
 OAI21_X1 _28267_ (.A(_09593_),
    .B1(_09585_),
    .B2(net420),
    .ZN(_02919_));
 NAND2_X1 _28268_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A2(_09584_),
    .ZN(_09594_));
 OAI21_X1 _28269_ (.A(_09594_),
    .B1(_09585_),
    .B2(_09498_),
    .ZN(_02920_));
 MUX2_X1 _28270_ (.A(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .B(net440),
    .S(_09582_),
    .Z(_02921_));
 MUX2_X1 _28271_ (.A(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .B(net333),
    .S(_09582_),
    .Z(_02922_));
 MUX2_X1 _28272_ (.A(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .B(net410),
    .S(_09582_),
    .Z(_02923_));
 NAND2_X1 _28273_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A2(_09584_),
    .ZN(_09595_));
 OAI21_X4 _28274_ (.A(_09595_),
    .B1(_09508_),
    .B2(_09585_),
    .ZN(_02924_));
 MUX2_X1 _28275_ (.A(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .B(_09445_),
    .S(_09582_),
    .Z(_02925_));
 NAND2_X1 _28276_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A2(_09584_),
    .ZN(_09596_));
 OAI21_X4 _28277_ (.A(_09596_),
    .B1(_09510_),
    .B2(_09585_),
    .ZN(_02926_));
 AND2_X1 _28278_ (.A1(_04604_),
    .A2(_09260_),
    .ZN(_09597_));
 BUF_X4 _28279_ (.A(_09597_),
    .Z(_09598_));
 BUF_X4 _28280_ (.A(_09598_),
    .Z(_09599_));
 MUX2_X1 _28281_ (.A(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .B(_05372_),
    .S(_09599_),
    .Z(_02927_));
 MUX2_X1 _28282_ (.A(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .B(_05410_),
    .S(_09599_),
    .Z(_02928_));
 NOR2_X1 _28283_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .A2(_05415_),
    .ZN(_09600_));
 AOI21_X1 _28284_ (.A(_09600_),
    .B1(_05850_),
    .B2(_05415_),
    .ZN(_02929_));
 NAND2_X2 _28285_ (.A1(_04604_),
    .A2(_09264_),
    .ZN(_09601_));
 CLKBUF_X3 _28286_ (.A(_09601_),
    .Z(_09602_));
 NAND2_X1 _28287_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .A2(_09602_),
    .ZN(_09603_));
 OAI21_X1 _28288_ (.A(_09603_),
    .B1(_09602_),
    .B2(_09475_),
    .ZN(_02930_));
 NAND2_X1 _28289_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .A2(_09602_),
    .ZN(_09604_));
 OAI21_X1 _28290_ (.A(_09604_),
    .B1(_09602_),
    .B2(_09477_),
    .ZN(_02931_));
 MUX2_X1 _28291_ (.A(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .B(_05544_),
    .S(_09599_),
    .Z(_02932_));
 MUX2_X1 _28292_ (.A(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .B(_05580_),
    .S(_09599_),
    .Z(_02933_));
 BUF_X4 _28293_ (.A(_09598_),
    .Z(_09605_));
 MUX2_X1 _28294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .B(_05614_),
    .S(_09605_),
    .Z(_02934_));
 MUX2_X1 _28295_ (.A(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .B(_05653_),
    .S(_09605_),
    .Z(_02935_));
 NOR2_X1 _28296_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .A2(_09599_),
    .ZN(_09606_));
 AOI21_X1 _28297_ (.A(_09606_),
    .B1(_09599_),
    .B2(_09384_),
    .ZN(_02936_));
 MUX2_X1 _28298_ (.A(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .B(_05721_),
    .S(_09605_),
    .Z(_02937_));
 MUX2_X1 _28299_ (.A(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .B(_05762_),
    .S(_09605_),
    .Z(_02938_));
 MUX2_X1 _28300_ (.A(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .B(_05802_),
    .S(_09605_),
    .Z(_02939_));
 MUX2_X1 _28301_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(_04855_),
    .Z(_02940_));
 NOR2_X1 _28302_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .A2(_09599_),
    .ZN(_09607_));
 AOI21_X1 _28303_ (.A(_09607_),
    .B1(_09599_),
    .B2(_06231_),
    .ZN(_02941_));
 MUX2_X1 _28304_ (.A(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .B(_05890_),
    .S(_09605_),
    .Z(_02942_));
 MUX2_X1 _28305_ (.A(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .B(_05928_),
    .S(_09605_),
    .Z(_02943_));
 MUX2_X1 _28306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .B(_09434_),
    .S(_09605_),
    .Z(_02944_));
 NOR2_X1 _28307_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .A2(_09599_),
    .ZN(_09608_));
 AOI21_X1 _28308_ (.A(_09608_),
    .B1(_09599_),
    .B2(_06234_),
    .ZN(_02945_));
 MUX2_X1 _28309_ (.A(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .B(_09438_),
    .S(_09605_),
    .Z(_02946_));
 MUX2_X1 _28310_ (.A(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .B(_09444_),
    .S(_09605_),
    .Z(_02947_));
 NAND2_X1 _28311_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .A2(_09602_),
    .ZN(_09609_));
 OAI21_X1 _28312_ (.A(_09609_),
    .B1(_09602_),
    .B2(_09484_),
    .ZN(_02948_));
 MUX2_X1 _28313_ (.A(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .B(_09460_),
    .S(_09598_),
    .Z(_02949_));
 MUX2_X1 _28314_ (.A(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .B(_09463_),
    .S(_09598_),
    .Z(_02950_));
 MUX2_X1 _28315_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(_04855_),
    .Z(_02951_));
 MUX2_X1 _28316_ (.A(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .B(_04602_),
    .S(_09598_),
    .Z(_02952_));
 MUX2_X1 _28317_ (.A(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .B(_09464_),
    .S(_09598_),
    .Z(_02953_));
 NAND2_X1 _28318_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .A2(_09601_),
    .ZN(_09610_));
 OAI21_X1 _28319_ (.A(_09610_),
    .B1(_09602_),
    .B2(net420),
    .ZN(_02954_));
 NAND2_X1 _28320_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .A2(_09601_),
    .ZN(_09611_));
 OAI21_X1 _28321_ (.A(_09611_),
    .B1(_09602_),
    .B2(_09498_),
    .ZN(_02955_));
 MUX2_X1 _28322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .B(_09467_),
    .S(_09598_),
    .Z(_02956_));
 MUX2_X1 _28323_ (.A(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .B(_04850_),
    .S(_09598_),
    .Z(_02957_));
 MUX2_X1 _28324_ (.A(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .B(_05094_),
    .S(_09598_),
    .Z(_02958_));
 NAND2_X1 _28325_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A2(_09601_),
    .ZN(_09612_));
 OAI21_X4 _28326_ (.A(_09612_),
    .B1(net447),
    .B2(_09602_),
    .ZN(_02959_));
 MUX2_X1 _28327_ (.A(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .B(_05211_),
    .S(_09598_),
    .Z(_02960_));
 NAND2_X1 _28328_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(_09601_),
    .ZN(_09613_));
 OAI21_X2 _28329_ (.A(_09613_),
    .B1(net438),
    .B2(_09602_),
    .ZN(_02961_));
 MUX2_X1 _28330_ (.A(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .B(_05974_),
    .S(_09558_),
    .Z(_02962_));
 MUX2_X1 _28331_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .S(_06246_),
    .Z(_02963_));
 AND2_X1 _28332_ (.A1(_05374_),
    .A2(_09260_),
    .ZN(_09614_));
 BUF_X4 _28333_ (.A(_09614_),
    .Z(_09615_));
 BUF_X4 _28334_ (.A(_09615_),
    .Z(_09616_));
 MUX2_X1 _28335_ (.A(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .B(_05372_),
    .S(_09616_),
    .Z(_02964_));
 MUX2_X1 _28336_ (.A(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .B(_05410_),
    .S(_09616_),
    .Z(_02965_));
 NAND2_X2 _28337_ (.A1(_05374_),
    .A2(_09264_),
    .ZN(_09617_));
 CLKBUF_X3 _28338_ (.A(_09617_),
    .Z(_09618_));
 NAND2_X1 _28339_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .A2(_09618_),
    .ZN(_09619_));
 OAI21_X1 _28340_ (.A(_09619_),
    .B1(_09618_),
    .B2(_09475_),
    .ZN(_02966_));
 NAND2_X1 _28341_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .A2(_09618_),
    .ZN(_09620_));
 OAI21_X1 _28342_ (.A(_09620_),
    .B1(_09618_),
    .B2(_09477_),
    .ZN(_02967_));
 MUX2_X1 _28343_ (.A(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .B(_05544_),
    .S(_09616_),
    .Z(_02968_));
 MUX2_X1 _28344_ (.A(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .B(_05580_),
    .S(_09616_),
    .Z(_02969_));
 BUF_X4 _28345_ (.A(_09615_),
    .Z(_09621_));
 MUX2_X1 _28346_ (.A(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .B(_05614_),
    .S(_09621_),
    .Z(_02970_));
 MUX2_X1 _28347_ (.A(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .B(_05653_),
    .S(_09621_),
    .Z(_02971_));
 NOR2_X1 _28348_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .A2(_09616_),
    .ZN(_09622_));
 AOI21_X1 _28349_ (.A(_09622_),
    .B1(_09616_),
    .B2(_06222_),
    .ZN(_02972_));
 MUX2_X1 _28350_ (.A(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .B(_05721_),
    .S(_09621_),
    .Z(_02973_));
 NOR2_X1 _28351_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .A2(_05415_),
    .ZN(_09623_));
 AOI21_X1 _28352_ (.A(_09623_),
    .B1(_06016_),
    .B2(_05415_),
    .ZN(_02974_));
 MUX2_X1 _28353_ (.A(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .B(_05762_),
    .S(_09621_),
    .Z(_02975_));
 MUX2_X1 _28354_ (.A(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .B(_05802_),
    .S(_09621_),
    .Z(_02976_));
 NOR2_X1 _28355_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .A2(_09616_),
    .ZN(_09624_));
 AOI21_X1 _28356_ (.A(_09624_),
    .B1(_09616_),
    .B2(_06231_),
    .ZN(_02977_));
 MUX2_X1 _28357_ (.A(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .B(_05890_),
    .S(_09621_),
    .Z(_02978_));
 MUX2_X1 _28358_ (.A(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .B(_05928_),
    .S(_09621_),
    .Z(_02979_));
 MUX2_X1 _28359_ (.A(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .B(_05974_),
    .S(_09621_),
    .Z(_02980_));
 NOR2_X1 _28360_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .A2(_09616_),
    .ZN(_09625_));
 AOI21_X1 _28361_ (.A(_09625_),
    .B1(_09616_),
    .B2(_06234_),
    .ZN(_02981_));
 MUX2_X1 _28362_ (.A(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .B(_06062_),
    .S(_09621_),
    .Z(_02982_));
 MUX2_X1 _28363_ (.A(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .B(_06100_),
    .S(_09621_),
    .Z(_02983_));
 NAND2_X1 _28364_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .A2(_09618_),
    .ZN(_09626_));
 OAI21_X1 _28365_ (.A(_09626_),
    .B1(_09618_),
    .B2(_09484_),
    .ZN(_02984_));
 MUX2_X1 _28366_ (.A(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .B(_06062_),
    .S(_09558_),
    .Z(_02985_));
 MUX2_X1 _28367_ (.A(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .B(_06174_),
    .S(_09615_),
    .Z(_02986_));
 MUX2_X1 _28368_ (.A(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .B(_06207_),
    .S(_09615_),
    .Z(_02987_));
 MUX2_X1 _28369_ (.A(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .B(_04602_),
    .S(_09615_),
    .Z(_02988_));
 MUX2_X1 _28370_ (.A(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .B(_04766_),
    .S(_09615_),
    .Z(_02989_));
 NAND2_X1 _28371_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .A2(_09617_),
    .ZN(_09627_));
 OAI21_X1 _28372_ (.A(_09627_),
    .B1(_09618_),
    .B2(_09488_),
    .ZN(_02990_));
 NAND2_X1 _28373_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .A2(_09617_),
    .ZN(_09628_));
 OAI21_X1 _28374_ (.A(_09628_),
    .B1(_09618_),
    .B2(_09498_),
    .ZN(_02991_));
 MUX2_X1 _28375_ (.A(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .B(_05037_),
    .S(_09615_),
    .Z(_02992_));
 MUX2_X1 _28376_ (.A(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .B(_04850_),
    .S(_09615_),
    .Z(_02993_));
 MUX2_X1 _28377_ (.A(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .B(_05094_),
    .S(_09615_),
    .Z(_02994_));
 NAND2_X1 _28378_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .A2(_09617_),
    .ZN(_09629_));
 OAI21_X4 _28379_ (.A(_09629_),
    .B1(_09508_),
    .B2(_09618_),
    .ZN(_02995_));
 MUX2_X1 _28380_ (.A(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .B(_06100_),
    .S(_09558_),
    .Z(_02996_));
 MUX2_X1 _28381_ (.A(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .B(net400),
    .S(_09615_),
    .Z(_02997_));
 NAND2_X1 _28382_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A2(_09617_),
    .ZN(_09630_));
 OAI21_X4 _28383_ (.A(_09630_),
    .B1(_09510_),
    .B2(_09618_),
    .ZN(_02998_));
 AND2_X1 _28384_ (.A1(_06214_),
    .A2(_09260_),
    .ZN(_09631_));
 BUF_X4 _28385_ (.A(_09631_),
    .Z(_09632_));
 BUF_X4 _28386_ (.A(_09632_),
    .Z(_09633_));
 MUX2_X1 _28387_ (.A(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .B(_05372_),
    .S(_09633_),
    .Z(_02999_));
 MUX2_X1 _28388_ (.A(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .B(_05410_),
    .S(_09633_),
    .Z(_03000_));
 NAND2_X2 _28389_ (.A1(_06214_),
    .A2(_09264_),
    .ZN(_09634_));
 CLKBUF_X3 _28390_ (.A(_09634_),
    .Z(_09635_));
 NAND2_X1 _28391_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .A2(_09635_),
    .ZN(_09636_));
 OAI21_X1 _28392_ (.A(_09636_),
    .B1(_09635_),
    .B2(_09475_),
    .ZN(_03001_));
 NAND2_X1 _28393_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .A2(_09635_),
    .ZN(_09637_));
 OAI21_X1 _28394_ (.A(_09637_),
    .B1(_09635_),
    .B2(_09477_),
    .ZN(_03002_));
 MUX2_X1 _28395_ (.A(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .B(_05544_),
    .S(_09633_),
    .Z(_03003_));
 MUX2_X1 _28396_ (.A(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .B(_05580_),
    .S(_09633_),
    .Z(_03004_));
 BUF_X4 _28397_ (.A(_09632_),
    .Z(_09638_));
 MUX2_X1 _28398_ (.A(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .B(_05614_),
    .S(_09638_),
    .Z(_03005_));
 MUX2_X1 _28399_ (.A(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .B(_05653_),
    .S(_09638_),
    .Z(_03006_));
 NAND2_X1 _28400_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .A2(_05803_),
    .ZN(_09639_));
 OAI21_X1 _28401_ (.A(_09639_),
    .B1(_06138_),
    .B2(_05806_),
    .ZN(_03007_));
 NOR2_X1 _28402_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .A2(_09633_),
    .ZN(_09640_));
 AOI21_X1 _28403_ (.A(_09640_),
    .B1(_09633_),
    .B2(_06222_),
    .ZN(_03008_));
 MUX2_X1 _28404_ (.A(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .B(_05721_),
    .S(_09638_),
    .Z(_03009_));
 MUX2_X1 _28405_ (.A(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .B(_05762_),
    .S(_09638_),
    .Z(_03010_));
 MUX2_X1 _28406_ (.A(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .B(_05802_),
    .S(_09638_),
    .Z(_03011_));
 NOR2_X1 _28407_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .A2(_09633_),
    .ZN(_09641_));
 AOI21_X1 _28408_ (.A(_09641_),
    .B1(_09633_),
    .B2(_06231_),
    .ZN(_03012_));
 MUX2_X1 _28409_ (.A(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .B(_05890_),
    .S(_09638_),
    .Z(_03013_));
 MUX2_X1 _28410_ (.A(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .B(_05928_),
    .S(_09638_),
    .Z(_03014_));
 MUX2_X1 _28411_ (.A(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .B(_05974_),
    .S(_09638_),
    .Z(_03015_));
 NOR2_X1 _28412_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .A2(_09633_),
    .ZN(_09642_));
 AOI21_X1 _28413_ (.A(_09642_),
    .B1(_09633_),
    .B2(_06234_),
    .ZN(_03016_));
 MUX2_X1 _28414_ (.A(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .B(_06062_),
    .S(_09638_),
    .Z(_03017_));
 MUX2_X1 _28415_ (.A(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .B(net405),
    .S(_09558_),
    .Z(_03018_));
 MUX2_X1 _28416_ (.A(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .B(_06100_),
    .S(_09638_),
    .Z(_03019_));
 NAND2_X1 _28417_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .A2(_09635_),
    .ZN(_09643_));
 OAI21_X1 _28418_ (.A(_09643_),
    .B1(_09635_),
    .B2(_09484_),
    .ZN(_03020_));
 MUX2_X1 _28419_ (.A(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .B(_06174_),
    .S(_09632_),
    .Z(_03021_));
 MUX2_X1 _28420_ (.A(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .B(_06207_),
    .S(_09632_),
    .Z(_03022_));
 MUX2_X1 _28421_ (.A(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .B(_04602_),
    .S(_09632_),
    .Z(_03023_));
 MUX2_X1 _28422_ (.A(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .B(_04766_),
    .S(_09632_),
    .Z(_03024_));
 NAND2_X1 _28423_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .A2(_09634_),
    .ZN(_09644_));
 OAI21_X1 _28424_ (.A(_09644_),
    .B1(_09635_),
    .B2(net420),
    .ZN(_03025_));
 NAND2_X1 _28425_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .A2(_09634_),
    .ZN(_09645_));
 OAI21_X1 _28426_ (.A(_09645_),
    .B1(_09635_),
    .B2(_09498_),
    .ZN(_03026_));
 MUX2_X1 _28427_ (.A(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .B(_05037_),
    .S(_09632_),
    .Z(_03027_));
 MUX2_X1 _28428_ (.A(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .B(net333),
    .S(_09632_),
    .Z(_03028_));
 MUX2_X1 _28429_ (.A(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .B(_06207_),
    .S(_09558_),
    .Z(_03029_));
 MUX2_X1 _28430_ (.A(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .B(_05094_),
    .S(_09632_),
    .Z(_03030_));
 NAND2_X1 _28431_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .A2(_09634_),
    .ZN(_09646_));
 OAI21_X4 _28432_ (.A(_09646_),
    .B1(_09508_),
    .B2(_09635_),
    .ZN(_03031_));
 MUX2_X1 _28433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .B(net400),
    .S(_09632_),
    .Z(_03032_));
 NAND2_X1 _28434_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .A2(_09634_),
    .ZN(_09647_));
 OAI21_X4 _28435_ (.A(_09647_),
    .B1(_09510_),
    .B2(_09635_),
    .ZN(_03033_));
 NAND2_X4 _28436_ (.A1(_04613_),
    .A2(_09420_),
    .ZN(_09648_));
 BUF_X4 _28437_ (.A(_09648_),
    .Z(_09649_));
 MUX2_X1 _28438_ (.A(_05372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .S(_09649_),
    .Z(_03034_));
 MUX2_X1 _28439_ (.A(_05410_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .S(_09649_),
    .Z(_03035_));
 BUF_X4 _28440_ (.A(_09648_),
    .Z(_09650_));
 NAND2_X1 _28441_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .A2(_09650_),
    .ZN(_09651_));
 BUF_X4 _28442_ (.A(_09648_),
    .Z(_09652_));
 OAI21_X1 _28443_ (.A(_09651_),
    .B1(_09652_),
    .B2(_05463_),
    .ZN(_03036_));
 NAND2_X1 _28444_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .A2(_09650_),
    .ZN(_09653_));
 OAI21_X1 _28445_ (.A(_09653_),
    .B1(_09652_),
    .B2(_05509_),
    .ZN(_03037_));
 MUX2_X1 _28446_ (.A(_05544_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .S(_09649_),
    .Z(_03038_));
 MUX2_X1 _28447_ (.A(_09370_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .S(_09649_),
    .Z(_03039_));
 MUX2_X1 _28448_ (.A(_09359_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(_04855_),
    .Z(_03040_));
 MUX2_X1 _28449_ (.A(_05614_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .S(_09649_),
    .Z(_03041_));
 MUX2_X1 _28450_ (.A(_09377_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .S(_09649_),
    .Z(_03042_));
 NAND2_X1 _28451_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .A2(_09650_),
    .ZN(_09654_));
 OAI21_X1 _28452_ (.A(_09654_),
    .B1(_09652_),
    .B2(_05687_),
    .ZN(_03043_));
 MUX2_X1 _28453_ (.A(_09372_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .S(_09649_),
    .Z(_03044_));
 MUX2_X1 _28454_ (.A(_05762_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .S(_09649_),
    .Z(_03045_));
 MUX2_X1 _28455_ (.A(_05802_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .S(_09649_),
    .Z(_03046_));
 NAND2_X1 _28456_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .A2(_09650_),
    .ZN(_09655_));
 OAI21_X1 _28457_ (.A(_09655_),
    .B1(_09652_),
    .B2(_05849_),
    .ZN(_03047_));
 MUX2_X1 _28458_ (.A(_09374_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .S(_09649_),
    .Z(_03048_));
 BUF_X4 _28459_ (.A(_09648_),
    .Z(_09656_));
 MUX2_X1 _28460_ (.A(_09375_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .S(_09656_),
    .Z(_03049_));
 MUX2_X1 _28461_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .S(_09656_),
    .Z(_03050_));
 MUX2_X1 _28462_ (.A(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .B(_04766_),
    .S(_09558_),
    .Z(_03051_));
 NAND2_X1 _28463_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .A2(_09650_),
    .ZN(_09657_));
 OAI21_X1 _28464_ (.A(_09657_),
    .B1(_09652_),
    .B2(_06015_),
    .ZN(_03052_));
 MUX2_X1 _28465_ (.A(_06062_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .S(_09656_),
    .Z(_03053_));
 MUX2_X1 _28466_ (.A(_06100_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .S(_09656_),
    .Z(_03054_));
 NAND2_X1 _28467_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .A2(_09650_),
    .ZN(_09658_));
 OAI21_X1 _28468_ (.A(_09658_),
    .B1(_09652_),
    .B2(_06137_),
    .ZN(_03055_));
 MUX2_X1 _28469_ (.A(net405),
    .B(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .S(_09656_),
    .Z(_03056_));
 MUX2_X1 _28470_ (.A(_06207_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .S(_09656_),
    .Z(_03057_));
 MUX2_X1 _28471_ (.A(_04601_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .S(_09656_),
    .Z(_03058_));
 MUX2_X1 _28472_ (.A(_04765_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .S(_09656_),
    .Z(_03059_));
 NAND2_X1 _28473_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A2(_09650_),
    .ZN(_09659_));
 OAI21_X1 _28474_ (.A(_09659_),
    .B1(_09652_),
    .B2(_04907_),
    .ZN(_03060_));
 NAND2_X1 _28475_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A2(_09650_),
    .ZN(_09660_));
 OAI21_X1 _28476_ (.A(_09660_),
    .B1(_09652_),
    .B2(_04977_),
    .ZN(_03061_));
 NAND2_X1 _28477_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .A2(_05803_),
    .ZN(_09661_));
 OAI21_X1 _28478_ (.A(_09661_),
    .B1(_04908_),
    .B2(_05806_),
    .ZN(_03062_));
 MUX2_X1 _28479_ (.A(_05036_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .S(_09656_),
    .Z(_03063_));
 MUX2_X1 _28480_ (.A(_04849_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .S(_09656_),
    .Z(_03064_));
 MUX2_X1 _28481_ (.A(_05093_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .S(_09648_),
    .Z(_03065_));
 NAND2_X1 _28482_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A2(_09650_),
    .ZN(_09662_));
 OAI21_X4 _28483_ (.A(_09662_),
    .B1(_05147_),
    .B2(_09652_),
    .ZN(_03066_));
 MUX2_X1 _28484_ (.A(_05210_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .S(_09648_),
    .Z(_03067_));
 NAND2_X1 _28485_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A2(_09650_),
    .ZN(_09663_));
 OAI21_X1 _28486_ (.A(_09663_),
    .B1(_09652_),
    .B2(_05259_),
    .ZN(_03068_));
 MUX2_X1 _28487_ (.A(_05371_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .S(_04615_),
    .Z(_03069_));
 MUX2_X1 _28488_ (.A(_05409_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .S(_04615_),
    .Z(_03070_));
 NAND2_X1 _28489_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .A2(_04856_),
    .ZN(_09664_));
 OAI21_X1 _28490_ (.A(_09664_),
    .B1(_05464_),
    .B2(_04909_),
    .ZN(_03071_));
 NAND2_X1 _28491_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .A2(_04856_),
    .ZN(_09665_));
 OAI21_X1 _28492_ (.A(_09665_),
    .B1(_05510_),
    .B2(_04909_),
    .ZN(_03072_));
 NAND2_X1 _28493_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .A2(_05803_),
    .ZN(_09666_));
 OAI21_X2 _28494_ (.A(_09666_),
    .B1(net442),
    .B2(_05803_),
    .ZN(_03073_));
 NOR2_X1 _28495_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .A2(_09177_),
    .ZN(_09667_));
 AOI21_X1 _28496_ (.A(_09667_),
    .B1(_09177_),
    .B2(_06222_),
    .ZN(_03074_));
 MUX2_X1 _28497_ (.A(_05543_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .S(_04615_),
    .Z(_03075_));
 MUX2_X1 _28498_ (.A(_05579_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .S(_04615_),
    .Z(_03076_));
 BUF_X4 _28499_ (.A(_04614_),
    .Z(_09668_));
 MUX2_X1 _28500_ (.A(_05613_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .S(_09668_),
    .Z(_03077_));
 MUX2_X1 _28501_ (.A(_05652_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .S(_09668_),
    .Z(_03078_));
 NAND2_X1 _28502_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .A2(_04856_),
    .ZN(_09669_));
 OAI21_X1 _28503_ (.A(_09669_),
    .B1(_05688_),
    .B2(_04909_),
    .ZN(_03079_));
 MUX2_X1 _28504_ (.A(_05720_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .S(_09668_),
    .Z(_03080_));
 MUX2_X1 _28505_ (.A(_05761_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .S(_09668_),
    .Z(_03081_));
 MUX2_X1 _28506_ (.A(_05801_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .S(_09668_),
    .Z(_03082_));
 NAND2_X1 _28507_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .A2(_04856_),
    .ZN(_09670_));
 OAI21_X1 _28508_ (.A(_09670_),
    .B1(_05850_),
    .B2(_04909_),
    .ZN(_03083_));
 MUX2_X1 _28509_ (.A(_05889_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .S(_09668_),
    .Z(_03084_));
 MUX2_X1 _28510_ (.A(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .B(_05037_),
    .S(_05414_),
    .Z(_03085_));
 MUX2_X1 _28511_ (.A(_05927_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .S(_09668_),
    .Z(_03086_));
 MUX2_X1 _28512_ (.A(_05973_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .S(_09668_),
    .Z(_03087_));
 NAND2_X1 _28513_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .A2(_04856_),
    .ZN(_09671_));
 OAI21_X1 _28514_ (.A(_09671_),
    .B1(_06016_),
    .B2(_04909_),
    .ZN(_03088_));
 MUX2_X1 _28515_ (.A(_06061_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .S(_09668_),
    .Z(_03089_));
 MUX2_X1 _28516_ (.A(_06099_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .S(_09668_),
    .Z(_03090_));
 NAND2_X1 _28517_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .A2(_04856_),
    .ZN(_09672_));
 OAI21_X1 _28518_ (.A(_09672_),
    .B1(_06138_),
    .B2(_04909_),
    .ZN(_03091_));
 MUX2_X1 _28519_ (.A(_06173_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .S(_04614_),
    .Z(_03092_));
 MUX2_X1 _28520_ (.A(_06206_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .S(_04614_),
    .Z(_01184_));
 MUX2_X1 _28521_ (.A(net107),
    .B(net122),
    .S(_03961_),
    .Z(_09673_));
 OR2_X1 _28522_ (.A1(_03978_),
    .A2(_09673_),
    .ZN(_09674_));
 MUX2_X1 _28523_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(_03962_),
    .Z(_09675_));
 OAI21_X4 _28524_ (.A(_09674_),
    .B1(_09675_),
    .B2(_03965_),
    .ZN(_09676_));
 MUX2_X1 _28525_ (.A(net108),
    .B(net123),
    .S(_03961_),
    .Z(_09677_));
 OR2_X1 _28526_ (.A1(_03973_),
    .A2(_09677_),
    .ZN(_09678_));
 MUX2_X1 _28527_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(_03961_),
    .Z(_09679_));
 OAI21_X2 _28528_ (.A(_09678_),
    .B1(_09679_),
    .B2(_03965_),
    .ZN(_09680_));
 BUF_X4 _28529_ (.A(_09680_),
    .Z(_09681_));
 BUF_X4 _28530_ (.A(\cs_registers_i.pc_if_i[1] ),
    .Z(_09682_));
 MUX2_X1 _28531_ (.A(net110),
    .B(net126),
    .S(_09682_),
    .Z(_09683_));
 OR2_X1 _28532_ (.A1(_03973_),
    .A2(_09683_),
    .ZN(_09684_));
 MUX2_X2 _28533_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(_09682_),
    .Z(_09685_));
 OAI21_X4 _28534_ (.A(_09684_),
    .B1(_09685_),
    .B2(_03965_),
    .ZN(_09686_));
 NAND2_X4 _28535_ (.A1(_09681_),
    .A2(_09686_),
    .ZN(_09687_));
 MUX2_X1 _28536_ (.A(net109),
    .B(net125),
    .S(_09682_),
    .Z(_09688_));
 MUX2_X1 _28537_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(_03961_),
    .Z(_09689_));
 MUX2_X1 _28538_ (.A(_09688_),
    .B(_09689_),
    .S(_03973_),
    .Z(_09690_));
 BUF_X4 _28539_ (.A(_09690_),
    .Z(_09691_));
 NOR2_X4 _28540_ (.A1(_09687_),
    .A2(_09691_),
    .ZN(_09692_));
 BUF_X4 _28541_ (.A(_09692_),
    .Z(_09693_));
 NAND2_X2 _28542_ (.A1(_09676_),
    .A2(_09693_),
    .ZN(_09694_));
 CLKBUF_X3 _28543_ (.A(_09681_),
    .Z(_09695_));
 MUX2_X2 _28544_ (.A(_09683_),
    .B(_09685_),
    .S(_03973_),
    .Z(_09696_));
 CLKBUF_X3 _28545_ (.A(_09696_),
    .Z(_09697_));
 BUF_X4 _28546_ (.A(_09691_),
    .Z(_09698_));
 BUF_X4 _28547_ (.A(_09698_),
    .Z(_09699_));
 MUX2_X1 _28548_ (.A(net132),
    .B(net118),
    .S(_03961_),
    .Z(_09700_));
 MUX2_X1 _28549_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(_03961_),
    .Z(_09701_));
 MUX2_X1 _28550_ (.A(_09700_),
    .B(_09701_),
    .S(_03978_),
    .Z(_09702_));
 BUF_X4 _28551_ (.A(_09702_),
    .Z(_09703_));
 INV_X1 _28552_ (.A(_09703_),
    .ZN(_09704_));
 MUX2_X1 _28553_ (.A(net133),
    .B(net119),
    .S(_09682_),
    .Z(_09705_));
 MUX2_X1 _28554_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(_03961_),
    .Z(_09706_));
 MUX2_X2 _28555_ (.A(_09705_),
    .B(_09706_),
    .S(_03973_),
    .Z(_09707_));
 MUX2_X1 _28556_ (.A(net131),
    .B(net117),
    .S(_09682_),
    .Z(_09708_));
 MUX2_X1 _28557_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(_09682_),
    .Z(_09709_));
 MUX2_X2 _28558_ (.A(_09708_),
    .B(_09709_),
    .S(_03964_),
    .Z(_09710_));
 MUX2_X1 _28559_ (.A(net106),
    .B(net121),
    .S(_09682_),
    .Z(_09711_));
 MUX2_X1 _28560_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(_09682_),
    .Z(_09712_));
 MUX2_X2 _28561_ (.A(_09711_),
    .B(_09712_),
    .S(_03973_),
    .Z(_09713_));
 MUX2_X1 _28562_ (.A(net105),
    .B(net120),
    .S(_09682_),
    .Z(_09714_));
 MUX2_X1 _28563_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(_09682_),
    .Z(_09715_));
 MUX2_X2 _28564_ (.A(_09714_),
    .B(_09715_),
    .S(_03973_),
    .Z(_09716_));
 NOR4_X4 _28565_ (.A1(_09707_),
    .A2(_09710_),
    .A3(_09713_),
    .A4(_09716_),
    .ZN(_09717_));
 NAND2_X1 _28566_ (.A1(_09704_),
    .A2(_09717_),
    .ZN(_09718_));
 BUF_X4 _28567_ (.A(_09686_),
    .Z(_09719_));
 MUX2_X1 _28568_ (.A(net130),
    .B(net116),
    .S(_03962_),
    .Z(_09720_));
 MUX2_X1 _28569_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(_03962_),
    .Z(_09721_));
 MUX2_X2 _28570_ (.A(_09720_),
    .B(_09721_),
    .S(_03978_),
    .Z(_09722_));
 MUX2_X1 _28571_ (.A(net129),
    .B(net115),
    .S(_03961_),
    .Z(_09723_));
 MUX2_X1 _28572_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(_03961_),
    .Z(_09724_));
 MUX2_X1 _28573_ (.A(_09723_),
    .B(_09724_),
    .S(_03978_),
    .Z(_09725_));
 CLKBUF_X3 _28574_ (.A(_09725_),
    .Z(_09726_));
 NOR2_X1 _28575_ (.A1(_09722_),
    .A2(_09726_),
    .ZN(_09727_));
 MUX2_X1 _28576_ (.A(net124),
    .B(net111),
    .S(_03962_),
    .Z(_09728_));
 MUX2_X1 _28577_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(_03962_),
    .Z(_09729_));
 MUX2_X1 _28578_ (.A(_09728_),
    .B(_09729_),
    .S(_03978_),
    .Z(_09730_));
 MUX2_X1 _28579_ (.A(net127),
    .B(net112),
    .S(_03962_),
    .Z(_09731_));
 MUX2_X1 _28580_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(_03962_),
    .Z(_09732_));
 MUX2_X2 _28581_ (.A(_09731_),
    .B(_09732_),
    .S(_03978_),
    .Z(_09733_));
 MUX2_X1 _28582_ (.A(net128),
    .B(net114),
    .S(_03962_),
    .Z(_09734_));
 MUX2_X1 _28583_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(_03962_),
    .Z(_09735_));
 MUX2_X1 _28584_ (.A(_09734_),
    .B(_09735_),
    .S(_03978_),
    .Z(_09736_));
 NOR3_X1 _28585_ (.A1(_09730_),
    .A2(_09733_),
    .A3(_09736_),
    .ZN(_09737_));
 NAND2_X1 _28586_ (.A1(_09727_),
    .A2(_09737_),
    .ZN(_09738_));
 NOR2_X1 _28587_ (.A1(_09691_),
    .A2(_09738_),
    .ZN(_09739_));
 AOI21_X1 _28588_ (.A(_09719_),
    .B1(_09676_),
    .B2(_09739_),
    .ZN(_09740_));
 OAI221_X1 _28589_ (.A(_09695_),
    .B1(_09697_),
    .B2(_09699_),
    .C1(_09718_),
    .C2(_09740_),
    .ZN(_09741_));
 MUX2_X1 _28590_ (.A(net104),
    .B(_03968_),
    .S(_03963_),
    .Z(_09742_));
 MUX2_X1 _28591_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(_03963_),
    .Z(_09743_));
 MUX2_X1 _28592_ (.A(_09742_),
    .B(_09743_),
    .S(_03979_),
    .Z(_09744_));
 BUF_X4 _28593_ (.A(_09744_),
    .Z(_09745_));
 MUX2_X1 _28594_ (.A(net113),
    .B(_03967_),
    .S(_03963_),
    .Z(_09746_));
 OR2_X1 _28595_ (.A1(_03979_),
    .A2(_09746_),
    .ZN(_09747_));
 MUX2_X1 _28596_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(_03963_),
    .Z(_09748_));
 BUF_X4 _28597_ (.A(_03965_),
    .Z(_09749_));
 OAI21_X4 _28598_ (.A(_09747_),
    .B1(_09748_),
    .B2(_09749_),
    .ZN(_09750_));
 NOR2_X1 _28599_ (.A1(_09745_),
    .A2(_09750_),
    .ZN(_09751_));
 CLKBUF_X3 _28600_ (.A(_09751_),
    .Z(_09752_));
 NAND3_X1 _28601_ (.A1(_09694_),
    .A2(_09741_),
    .A3(_09752_),
    .ZN(_09753_));
 MUX2_X1 _28602_ (.A(_09673_),
    .B(_09675_),
    .S(_03979_),
    .Z(_09754_));
 CLKBUF_X3 _28603_ (.A(_09754_),
    .Z(_09755_));
 CLKBUF_X3 _28604_ (.A(_09755_),
    .Z(_09756_));
 NAND2_X2 _28605_ (.A1(_09686_),
    .A2(_09690_),
    .ZN(_09757_));
 NOR4_X1 _28606_ (.A1(_09695_),
    .A2(_09756_),
    .A3(_09738_),
    .A4(_09757_),
    .ZN(_09758_));
 NOR2_X1 _28607_ (.A1(_09686_),
    .A2(_09691_),
    .ZN(_09759_));
 NAND2_X2 _28608_ (.A1(_09681_),
    .A2(_09759_),
    .ZN(_09760_));
 OR2_X1 _28609_ (.A1(_07136_),
    .A2(_09714_),
    .ZN(_09761_));
 OAI21_X4 _28610_ (.A(_09761_),
    .B1(_09715_),
    .B2(_09749_),
    .ZN(_09762_));
 CLKBUF_X3 _28611_ (.A(_09713_),
    .Z(_09763_));
 AOI21_X1 _28612_ (.A(_09760_),
    .B1(_09762_),
    .B2(_09763_),
    .ZN(_09764_));
 AOI21_X1 _28613_ (.A(_09758_),
    .B1(_09764_),
    .B2(_09756_),
    .ZN(_09765_));
 NAND2_X4 _28614_ (.A1(_09745_),
    .A2(_09750_),
    .ZN(_09766_));
 OR2_X1 _28615_ (.A1(_03979_),
    .A2(_09742_),
    .ZN(_09767_));
 OAI21_X4 _28616_ (.A(_09767_),
    .B1(_09743_),
    .B2(_03965_),
    .ZN(_09768_));
 NAND2_X4 _28617_ (.A1(_09768_),
    .A2(_09750_),
    .ZN(_09769_));
 MUX2_X2 _28618_ (.A(_09677_),
    .B(_09679_),
    .S(_03978_),
    .Z(_09770_));
 NOR2_X4 _28619_ (.A1(_09770_),
    .A2(_09696_),
    .ZN(_09771_));
 BUF_X4 _28620_ (.A(_09770_),
    .Z(_09772_));
 OR2_X1 _28621_ (.A1(_03973_),
    .A2(_09688_),
    .ZN(_09773_));
 OAI21_X4 _28622_ (.A(_09773_),
    .B1(_09689_),
    .B2(_03965_),
    .ZN(_09774_));
 BUF_X4 _28623_ (.A(_09774_),
    .Z(_09775_));
 NOR2_X4 _28624_ (.A1(_09772_),
    .A2(_09775_),
    .ZN(_09776_));
 NOR2_X4 _28625_ (.A1(_09771_),
    .A2(_09776_),
    .ZN(_09777_));
 BUF_X4 _28626_ (.A(_09777_),
    .Z(_09778_));
 INV_X1 _28627_ (.A(_09727_),
    .ZN(_09779_));
 NOR3_X1 _28628_ (.A1(_09779_),
    .A2(_09718_),
    .A3(_09694_),
    .ZN(_09780_));
 NOR2_X1 _28629_ (.A1(_09778_),
    .A2(_09780_),
    .ZN(_09781_));
 OAI221_X1 _28630_ (.A(_09753_),
    .B1(_09765_),
    .B2(_09766_),
    .C1(_09769_),
    .C2(_09781_),
    .ZN(_09782_));
 MUX2_X1 _28631_ (.A(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .B(_09782_),
    .S(_07218_),
    .Z(_01532_));
 BUF_X4 _28632_ (.A(_07240_),
    .Z(_09783_));
 NAND2_X1 _28633_ (.A1(_11419_),
    .A2(_09783_),
    .ZN(_09784_));
 INV_X1 _28634_ (.A(_03966_),
    .ZN(_09785_));
 NOR3_X1 _28635_ (.A1(_07137_),
    .A2(_03981_),
    .A3(_09785_),
    .ZN(_09786_));
 OAI21_X1 _28636_ (.A(_03966_),
    .B1(_00136_),
    .B2(_03974_),
    .ZN(_09787_));
 OR2_X1 _28637_ (.A1(_04158_),
    .A2(_09787_),
    .ZN(_09788_));
 AOI21_X1 _28638_ (.A(_03971_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B2(_03974_),
    .ZN(_09789_));
 OAI21_X1 _28639_ (.A(_09788_),
    .B1(_09789_),
    .B2(_07138_),
    .ZN(_09790_));
 AOI221_X2 _28640_ (.A(_09786_),
    .B1(_09790_),
    .B2(_03981_),
    .C1(_07137_),
    .C2(_03971_),
    .ZN(_09791_));
 OAI21_X1 _28641_ (.A(_09784_),
    .B1(_09791_),
    .B2(_09783_),
    .ZN(_01533_));
 NOR3_X1 _28642_ (.A1(_09749_),
    .A2(_07133_),
    .A3(_09785_),
    .ZN(_09792_));
 AOI21_X1 _28643_ (.A(_09792_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B2(_07133_),
    .ZN(_09793_));
 NOR3_X1 _28644_ (.A1(_07170_),
    .A2(_03971_),
    .A3(_09793_),
    .ZN(_09794_));
 MUX2_X1 _28645_ (.A(_08803_),
    .B(_09794_),
    .S(_07218_),
    .Z(_01534_));
 CLKBUF_X3 _28646_ (.A(_09745_),
    .Z(_09795_));
 MUX2_X2 _28647_ (.A(_09746_),
    .B(_09748_),
    .S(_03979_),
    .Z(_09796_));
 CLKBUF_X3 _28648_ (.A(_09796_),
    .Z(_09797_));
 CLKBUF_X3 _28649_ (.A(_09797_),
    .Z(_09798_));
 NAND2_X1 _28650_ (.A1(_09795_),
    .A2(_09798_),
    .ZN(_09799_));
 MUX2_X1 _28651_ (.A(_08813_),
    .B(_09799_),
    .S(_07218_),
    .Z(_01535_));
 CLKBUF_X3 _28652_ (.A(_09768_),
    .Z(_09800_));
 NAND2_X2 _28653_ (.A1(_09696_),
    .A2(_09774_),
    .ZN(_09801_));
 OAI21_X1 _28654_ (.A(_09695_),
    .B1(_09801_),
    .B2(_09797_),
    .ZN(_09802_));
 NAND2_X1 _28655_ (.A1(_09800_),
    .A2(_09802_),
    .ZN(_09803_));
 MUX2_X1 _28656_ (.A(_10291_),
    .B(_09803_),
    .S(_07218_),
    .Z(_01536_));
 MUX2_X1 _28657_ (.A(_09697_),
    .B(_09801_),
    .S(_09795_),
    .Z(_09804_));
 CLKBUF_X3 _28658_ (.A(_09716_),
    .Z(_09805_));
 OAI21_X1 _28659_ (.A(_09805_),
    .B1(_09766_),
    .B2(_09699_),
    .ZN(_09806_));
 BUF_X4 _28660_ (.A(_09772_),
    .Z(_09807_));
 CLKBUF_X3 _28661_ (.A(_09807_),
    .Z(_09808_));
 NOR2_X2 _28662_ (.A1(_09745_),
    .A2(_09772_),
    .ZN(_09809_));
 NAND2_X1 _28663_ (.A1(_09739_),
    .A2(_09809_),
    .ZN(_09810_));
 CLKBUF_X3 _28664_ (.A(_09719_),
    .Z(_09811_));
 OAI21_X1 _28665_ (.A(_09805_),
    .B1(_09810_),
    .B2(_09811_),
    .ZN(_09812_));
 AOI222_X2 _28666_ (.A1(_09762_),
    .A2(_09804_),
    .B1(_09806_),
    .B2(_09808_),
    .C1(_09798_),
    .C2(_09812_),
    .ZN(_09813_));
 MUX2_X1 _28667_ (.A(_10899_),
    .B(_09813_),
    .S(_07218_),
    .Z(_01537_));
 NAND2_X2 _28668_ (.A1(_09771_),
    .A2(_09775_),
    .ZN(_09814_));
 NOR2_X1 _28669_ (.A1(_09763_),
    .A2(_09814_),
    .ZN(_09815_));
 NOR2_X4 _28670_ (.A1(_09768_),
    .A2(_09796_),
    .ZN(_09816_));
 BUF_X4 _28671_ (.A(_09816_),
    .Z(_09817_));
 NOR2_X4 _28672_ (.A1(_09770_),
    .A2(_09801_),
    .ZN(_09818_));
 NAND2_X2 _28673_ (.A1(_09713_),
    .A2(_09716_),
    .ZN(_09819_));
 NOR2_X4 _28674_ (.A1(_09676_),
    .A2(_09819_),
    .ZN(_09820_));
 AND2_X2 _28675_ (.A1(_09818_),
    .A2(_09820_),
    .ZN(_09821_));
 OAI21_X1 _28676_ (.A(_09817_),
    .B1(_09821_),
    .B2(_09693_),
    .ZN(_09822_));
 CLKBUF_X3 _28677_ (.A(_09775_),
    .Z(_09823_));
 OAI21_X1 _28678_ (.A(_09752_),
    .B1(_09763_),
    .B2(_09823_),
    .ZN(_09824_));
 OAI21_X1 _28679_ (.A(_09822_),
    .B1(_09824_),
    .B2(_09687_),
    .ZN(_09825_));
 NOR2_X1 _28680_ (.A1(_09745_),
    .A2(_09687_),
    .ZN(_09826_));
 AOI21_X1 _28681_ (.A(_09826_),
    .B1(_09823_),
    .B2(_09745_),
    .ZN(_09827_));
 CLKBUF_X3 _28682_ (.A(_09750_),
    .Z(_09828_));
 MUX2_X1 _28683_ (.A(_09810_),
    .B(_09827_),
    .S(_09828_),
    .Z(_09829_));
 AOI21_X1 _28684_ (.A(_09825_),
    .B1(_09829_),
    .B2(_09763_),
    .ZN(_09830_));
 OR3_X1 _28685_ (.A1(_07253_),
    .A2(_09815_),
    .A3(_09830_),
    .ZN(_09831_));
 OAI21_X1 _28686_ (.A(_09831_),
    .B1(_07218_),
    .B2(_11062_),
    .ZN(_01538_));
 NAND2_X2 _28687_ (.A1(_09814_),
    .A2(_09816_),
    .ZN(_09832_));
 AOI21_X1 _28688_ (.A(_09819_),
    .B1(_09726_),
    .B2(_09722_),
    .ZN(_09833_));
 INV_X1 _28689_ (.A(_09833_),
    .ZN(_09834_));
 NOR2_X2 _28690_ (.A1(_09772_),
    .A2(_09686_),
    .ZN(_09835_));
 AOI22_X1 _28691_ (.A1(_09687_),
    .A2(_09755_),
    .B1(_09834_),
    .B2(_09835_),
    .ZN(_09836_));
 NOR2_X1 _28692_ (.A1(_09698_),
    .A2(_09836_),
    .ZN(_09837_));
 NOR2_X4 _28693_ (.A1(_09680_),
    .A2(_09757_),
    .ZN(_09838_));
 NAND2_X4 _28694_ (.A1(_09703_),
    .A2(_09717_),
    .ZN(_09839_));
 AND2_X2 _28695_ (.A1(_09838_),
    .A2(_09839_),
    .ZN(_09840_));
 CLKBUF_X3 _28696_ (.A(_09730_),
    .Z(_09841_));
 NOR2_X4 _28697_ (.A1(_09719_),
    .A2(_09775_),
    .ZN(_09842_));
 AOI221_X2 _28698_ (.A(_09837_),
    .B1(_09840_),
    .B2(_09841_),
    .C1(_09807_),
    .C2(_09842_),
    .ZN(_09843_));
 AOI22_X2 _28699_ (.A1(_09795_),
    .A2(_09756_),
    .B1(_09826_),
    .B2(_09823_),
    .ZN(_09844_));
 OAI222_X2 _28700_ (.A1(_09676_),
    .A2(_09803_),
    .B1(_09832_),
    .B2(_09843_),
    .C1(_09844_),
    .C2(_09828_),
    .ZN(_09845_));
 MUX2_X1 _28701_ (.A(_10477_),
    .B(_09845_),
    .S(_07218_),
    .Z(_01539_));
 OAI21_X1 _28702_ (.A(_09695_),
    .B1(_09823_),
    .B2(_09795_),
    .ZN(_09846_));
 NAND2_X1 _28703_ (.A1(_09766_),
    .A2(_09846_),
    .ZN(_09847_));
 NOR2_X4 _28704_ (.A1(_09681_),
    .A2(_09691_),
    .ZN(_09848_));
 NAND2_X1 _28705_ (.A1(_09755_),
    .A2(_09848_),
    .ZN(_09849_));
 INV_X1 _28706_ (.A(_09849_),
    .ZN(_09850_));
 AND2_X1 _28707_ (.A1(_09713_),
    .A2(_09818_),
    .ZN(_09851_));
 OR2_X1 _28708_ (.A1(_07136_),
    .A2(_09720_),
    .ZN(_09852_));
 OAI21_X4 _28709_ (.A(_09852_),
    .B1(_09721_),
    .B2(_09749_),
    .ZN(_09853_));
 OAI21_X1 _28710_ (.A(_09805_),
    .B1(_09755_),
    .B2(_09853_),
    .ZN(_09854_));
 AOI221_X2 _28711_ (.A(_09850_),
    .B1(_09851_),
    .B2(_09854_),
    .C1(_09840_),
    .C2(_09733_),
    .ZN(_09855_));
 OAI21_X1 _28712_ (.A(_09847_),
    .B1(_09855_),
    .B2(_09766_),
    .ZN(_09856_));
 MUX2_X1 _28713_ (.A(_10488_),
    .B(_09856_),
    .S(_07218_),
    .Z(_01540_));
 AOI21_X1 _28714_ (.A(_09699_),
    .B1(_09687_),
    .B2(_09828_),
    .ZN(_09857_));
 AOI21_X1 _28715_ (.A(_09795_),
    .B1(_09808_),
    .B2(_09699_),
    .ZN(_09858_));
 NAND2_X1 _28716_ (.A1(_09816_),
    .A2(_09849_),
    .ZN(_09859_));
 CLKBUF_X3 _28717_ (.A(_09736_),
    .Z(_09860_));
 AND2_X1 _28718_ (.A1(_09763_),
    .A2(_09805_),
    .ZN(_09861_));
 OAI21_X1 _28719_ (.A(_09861_),
    .B1(_09756_),
    .B2(_09727_),
    .ZN(_09862_));
 AOI221_X2 _28720_ (.A(_09859_),
    .B1(_09840_),
    .B2(_09860_),
    .C1(_09818_),
    .C2(_09862_),
    .ZN(_09863_));
 NOR3_X1 _28721_ (.A1(_09857_),
    .A2(_09858_),
    .A3(_09863_),
    .ZN(_09864_));
 BUF_X4 _28722_ (.A(_07180_),
    .Z(_09865_));
 MUX2_X1 _28723_ (.A(_10495_),
    .B(_09864_),
    .S(_09865_),
    .Z(_01541_));
 NAND2_X1 _28724_ (.A1(_10597_),
    .A2(_07253_),
    .ZN(_09866_));
 INV_X1 _28725_ (.A(_09710_),
    .ZN(_09867_));
 NAND2_X2 _28726_ (.A1(_09818_),
    .A2(_09820_),
    .ZN(_09868_));
 NAND2_X1 _28727_ (.A1(_09676_),
    .A2(_09738_),
    .ZN(_09869_));
 AOI21_X1 _28728_ (.A(_09719_),
    .B1(_09710_),
    .B2(_09869_),
    .ZN(_09870_));
 OAI21_X1 _28729_ (.A(_09681_),
    .B1(_09691_),
    .B2(_09870_),
    .ZN(_09871_));
 NOR2_X1 _28730_ (.A1(_09681_),
    .A2(_09696_),
    .ZN(_09872_));
 INV_X1 _28731_ (.A(_09872_),
    .ZN(_09873_));
 NAND3_X1 _28732_ (.A1(_09751_),
    .A2(_09871_),
    .A3(_09873_),
    .ZN(_09874_));
 NAND2_X1 _28733_ (.A1(_09726_),
    .A2(_09840_),
    .ZN(_09875_));
 NOR2_X1 _28734_ (.A1(_09692_),
    .A2(_09850_),
    .ZN(_09876_));
 NAND4_X1 _28735_ (.A1(_09868_),
    .A2(_09874_),
    .A3(_09875_),
    .A4(_09876_),
    .ZN(_09877_));
 NAND2_X1 _28736_ (.A1(_09814_),
    .A2(_09877_),
    .ZN(_09878_));
 NAND3_X1 _28737_ (.A1(_09868_),
    .A2(_09875_),
    .A3(_09876_),
    .ZN(_09879_));
 OAI22_X4 _28738_ (.A1(_09719_),
    .A2(_09774_),
    .B1(_09760_),
    .B2(_09820_),
    .ZN(_09880_));
 OAI21_X1 _28739_ (.A(_09817_),
    .B1(_09879_),
    .B2(_09880_),
    .ZN(_09881_));
 AOI22_X2 _28740_ (.A1(_09867_),
    .A2(_09878_),
    .B1(_09881_),
    .B2(_09874_),
    .ZN(_09882_));
 MUX2_X1 _28741_ (.A(_09697_),
    .B(_09710_),
    .S(_09776_),
    .Z(_09883_));
 NOR2_X4 _28742_ (.A1(_09745_),
    .A2(_09796_),
    .ZN(_09884_));
 NOR2_X1 _28743_ (.A1(_09828_),
    .A2(_09811_),
    .ZN(_09885_));
 AOI221_X2 _28744_ (.A(_09882_),
    .B1(_09883_),
    .B2(_09884_),
    .C1(_09795_),
    .C2(_09885_),
    .ZN(_09886_));
 OAI21_X1 _28745_ (.A(_09866_),
    .B1(_09886_),
    .B2(_09783_),
    .ZN(_01542_));
 BUF_X4 _28746_ (.A(_09884_),
    .Z(_09887_));
 NAND2_X2 _28747_ (.A1(_09695_),
    .A2(_09698_),
    .ZN(_09888_));
 MUX2_X1 _28748_ (.A(_03968_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(_03979_),
    .Z(_09889_));
 MUX2_X2 _28749_ (.A(_07334_),
    .B(_09889_),
    .S(_07169_),
    .Z(_09890_));
 NAND2_X2 _28750_ (.A1(_09687_),
    .A2(_09888_),
    .ZN(_09891_));
 OAI221_X2 _28751_ (.A(_09887_),
    .B1(_09888_),
    .B2(_09703_),
    .C1(_09890_),
    .C2(_09891_),
    .ZN(_09892_));
 AOI21_X1 _28752_ (.A(_09760_),
    .B1(_09869_),
    .B2(_09703_),
    .ZN(_09893_));
 OAI21_X1 _28753_ (.A(_09751_),
    .B1(_09890_),
    .B2(_09681_),
    .ZN(_09894_));
 NOR2_X1 _28754_ (.A1(_09893_),
    .A2(_09894_),
    .ZN(_09895_));
 NAND2_X1 _28755_ (.A1(_09816_),
    .A2(_09838_),
    .ZN(_09896_));
 AOI21_X1 _28756_ (.A(_09896_),
    .B1(_09839_),
    .B2(_09853_),
    .ZN(_09897_));
 NOR2_X1 _28757_ (.A1(_09895_),
    .A2(_09897_),
    .ZN(_09898_));
 AOI221_X2 _28758_ (.A(_09692_),
    .B1(_09821_),
    .B2(_09890_),
    .C1(_09848_),
    .C2(_09754_),
    .ZN(_09899_));
 INV_X1 _28759_ (.A(_09899_),
    .ZN(_09900_));
 OAI21_X1 _28760_ (.A(_09816_),
    .B1(_09880_),
    .B2(_09900_),
    .ZN(_09901_));
 NAND2_X1 _28761_ (.A1(_09898_),
    .A2(_09901_),
    .ZN(_09902_));
 AOI21_X1 _28762_ (.A(_09693_),
    .B1(_09898_),
    .B2(_09899_),
    .ZN(_09903_));
 OAI21_X1 _28763_ (.A(_09902_),
    .B1(_09903_),
    .B2(_09703_),
    .ZN(_09904_));
 NAND2_X1 _28764_ (.A1(_09797_),
    .A2(_09890_),
    .ZN(_09905_));
 AND2_X1 _28765_ (.A1(_09904_),
    .A2(_09905_),
    .ZN(_09906_));
 OAI221_X2 _28766_ (.A(_09892_),
    .B1(_09904_),
    .B2(_09828_),
    .C1(_09800_),
    .C2(_09906_),
    .ZN(_09907_));
 MUX2_X1 _28767_ (.A(_10759_),
    .B(_09907_),
    .S(_09865_),
    .Z(_01543_));
 NOR2_X1 _28768_ (.A1(_09840_),
    .A2(_09848_),
    .ZN(_09908_));
 NOR2_X1 _28769_ (.A1(_09676_),
    .A2(_09908_),
    .ZN(_09909_));
 NOR2_X2 _28770_ (.A1(_09692_),
    .A2(_09909_),
    .ZN(_09910_));
 MUX2_X1 _28771_ (.A(_03967_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(_03979_),
    .Z(_09911_));
 MUX2_X2 _28772_ (.A(_07346_),
    .B(_09911_),
    .S(_07169_),
    .Z(_09912_));
 AOI22_X2 _28773_ (.A1(_09707_),
    .A2(_09880_),
    .B1(_09912_),
    .B2(_09821_),
    .ZN(_09913_));
 AOI21_X2 _28774_ (.A(_09766_),
    .B1(_09910_),
    .B2(_09913_),
    .ZN(_09914_));
 NAND2_X1 _28775_ (.A1(_09768_),
    .A2(_09797_),
    .ZN(_09915_));
 NAND2_X1 _28776_ (.A1(_09807_),
    .A2(_09912_),
    .ZN(_09916_));
 AOI21_X1 _28777_ (.A(_09692_),
    .B1(_09818_),
    .B2(_09869_),
    .ZN(_09917_));
 AOI21_X1 _28778_ (.A(_09915_),
    .B1(_09916_),
    .B2(_09917_),
    .ZN(_09918_));
 AOI21_X1 _28779_ (.A(_09914_),
    .B1(_09912_),
    .B2(_09807_),
    .ZN(_09919_));
 NOR2_X1 _28780_ (.A1(_09693_),
    .A2(_09919_),
    .ZN(_09920_));
 OAI22_X2 _28781_ (.A1(_09914_),
    .A2(_09918_),
    .B1(_09920_),
    .B2(_09707_),
    .ZN(_09921_));
 AOI22_X2 _28782_ (.A1(_09776_),
    .A2(_09707_),
    .B1(_09912_),
    .B2(_09778_),
    .ZN(_09922_));
 INV_X1 _28783_ (.A(_09912_),
    .ZN(_09923_));
 OAI221_X2 _28784_ (.A(_09921_),
    .B1(_09922_),
    .B2(_09769_),
    .C1(_09799_),
    .C2(_09923_),
    .ZN(_09924_));
 MUX2_X1 _28785_ (.A(_10752_),
    .B(_09924_),
    .S(_09865_),
    .Z(_01544_));
 NAND2_X1 _28786_ (.A1(_10767_),
    .A2(_07253_),
    .ZN(_09925_));
 NAND2_X1 _28787_ (.A1(_07136_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .ZN(_09926_));
 NAND2_X1 _28788_ (.A1(_09749_),
    .A2(net111),
    .ZN(_09927_));
 AOI21_X1 _28789_ (.A(_03963_),
    .B1(_09926_),
    .B2(_09927_),
    .ZN(_09928_));
 AOI21_X2 _28790_ (.A(_09928_),
    .B1(_07358_),
    .B2(_03963_),
    .ZN(_09929_));
 OAI22_X1 _28791_ (.A1(_09762_),
    .A2(_09917_),
    .B1(_09929_),
    .B2(_09681_),
    .ZN(_09930_));
 AND2_X1 _28792_ (.A1(_09752_),
    .A2(_09930_),
    .ZN(_09931_));
 AOI21_X1 _28793_ (.A(_09772_),
    .B1(_09820_),
    .B2(_09929_),
    .ZN(_09932_));
 OAI21_X1 _28794_ (.A(_09696_),
    .B1(_09691_),
    .B2(_09932_),
    .ZN(_09933_));
 AOI21_X1 _28795_ (.A(_09797_),
    .B1(_09910_),
    .B2(_09933_),
    .ZN(_09934_));
 OAI22_X1 _28796_ (.A1(_09805_),
    .A2(_09814_),
    .B1(_09931_),
    .B2(_09934_),
    .ZN(_09935_));
 OAI21_X1 _28797_ (.A(_09935_),
    .B1(_09929_),
    .B2(_09828_),
    .ZN(_09936_));
 OAI21_X1 _28798_ (.A(_09888_),
    .B1(_09929_),
    .B2(_09771_),
    .ZN(_09937_));
 AOI221_X2 _28799_ (.A(_09931_),
    .B1(_09936_),
    .B2(_09795_),
    .C1(_09937_),
    .C2(_09887_),
    .ZN(_09938_));
 OAI21_X1 _28800_ (.A(_09925_),
    .B1(_09938_),
    .B2(_09783_),
    .ZN(_01545_));
 NAND2_X1 _28801_ (.A1(_07137_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .ZN(_09939_));
 NAND2_X1 _28802_ (.A1(_09749_),
    .A2(net112),
    .ZN(_09940_));
 NAND3_X1 _28803_ (.A1(_07170_),
    .A2(_09939_),
    .A3(_09940_),
    .ZN(_09941_));
 OAI21_X2 _28804_ (.A(_09941_),
    .B1(_07369_),
    .B2(_07170_),
    .ZN(_09942_));
 NOR2_X1 _28805_ (.A1(_09800_),
    .A2(_09828_),
    .ZN(_09943_));
 AOI21_X1 _28806_ (.A(_09943_),
    .B1(_09778_),
    .B2(_09887_),
    .ZN(_09944_));
 NAND2_X1 _28807_ (.A1(_09851_),
    .A2(_09869_),
    .ZN(_09945_));
 OAI221_X2 _28808_ (.A(_09945_),
    .B1(_09699_),
    .B2(_09687_),
    .C1(_09695_),
    .C2(_09942_),
    .ZN(_09946_));
 OAI21_X1 _28809_ (.A(_09910_),
    .B1(_09942_),
    .B2(_09868_),
    .ZN(_09947_));
 AOI22_X2 _28810_ (.A1(_09752_),
    .A2(_09946_),
    .B1(_09947_),
    .B2(_09817_),
    .ZN(_09948_));
 OAI22_X2 _28811_ (.A1(_09942_),
    .A2(_09944_),
    .B1(_09948_),
    .B2(_09815_),
    .ZN(_09949_));
 MUX2_X1 _28812_ (.A(_10750_),
    .B(_09949_),
    .S(_09865_),
    .Z(_01546_));
 NOR2_X1 _28813_ (.A1(_09766_),
    .A2(_09868_),
    .ZN(_09950_));
 AOI21_X1 _28814_ (.A(_09950_),
    .B1(_09778_),
    .B2(_09887_),
    .ZN(_09951_));
 MUX2_X1 _28815_ (.A(_10290_),
    .B(_09951_),
    .S(_09865_),
    .Z(_01547_));
 NAND2_X1 _28816_ (.A1(_11935_),
    .A2(_07253_),
    .ZN(_09952_));
 MUX2_X1 _28817_ (.A(net114),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(_03979_),
    .Z(_09953_));
 MUX2_X2 _28818_ (.A(_07382_),
    .B(_09953_),
    .S(_07169_),
    .Z(_09954_));
 NAND2_X1 _28819_ (.A1(_09772_),
    .A2(_09954_),
    .ZN(_09955_));
 AND2_X1 _28820_ (.A1(_09727_),
    .A2(_09737_),
    .ZN(_09956_));
 NAND3_X1 _28821_ (.A1(_09755_),
    .A2(_09818_),
    .A3(_09956_),
    .ZN(_09957_));
 OAI21_X1 _28822_ (.A(_09681_),
    .B1(_09719_),
    .B2(_09841_),
    .ZN(_09958_));
 NOR2_X1 _28823_ (.A1(_09696_),
    .A2(_09775_),
    .ZN(_09959_));
 OAI221_X1 _28824_ (.A(_09955_),
    .B1(_09957_),
    .B2(_09718_),
    .C1(_09958_),
    .C2(_09959_),
    .ZN(_09960_));
 MUX2_X1 _28825_ (.A(_09841_),
    .B(_09954_),
    .S(_09820_),
    .Z(_09961_));
 AOI22_X1 _28826_ (.A1(_09841_),
    .A2(_09959_),
    .B1(_09961_),
    .B2(_09759_),
    .ZN(_09962_));
 OAI21_X1 _28827_ (.A(_09910_),
    .B1(_09962_),
    .B2(_09807_),
    .ZN(_09963_));
 AOI22_X1 _28828_ (.A1(_09752_),
    .A2(_09960_),
    .B1(_09963_),
    .B2(_09817_),
    .ZN(_09964_));
 INV_X1 _28829_ (.A(_09841_),
    .ZN(_09965_));
 AOI21_X1 _28830_ (.A(_09964_),
    .B1(_09965_),
    .B2(_09693_),
    .ZN(_09966_));
 AOI22_X1 _28831_ (.A1(_09776_),
    .A2(_09841_),
    .B1(_09954_),
    .B2(_09823_),
    .ZN(_09967_));
 OAI21_X1 _28832_ (.A(_09955_),
    .B1(_09967_),
    .B2(_09811_),
    .ZN(_09968_));
 AOI221_X2 _28833_ (.A(_09966_),
    .B1(_09954_),
    .B2(_09943_),
    .C1(_09887_),
    .C2(_09968_),
    .ZN(_09969_));
 OAI21_X1 _28834_ (.A(_09952_),
    .B1(_09969_),
    .B2(_09783_),
    .ZN(_01548_));
 AND2_X1 _28835_ (.A1(_09755_),
    .A2(_09840_),
    .ZN(_09970_));
 OR2_X1 _28836_ (.A1(_07136_),
    .A2(_09731_),
    .ZN(_09971_));
 OAI21_X2 _28837_ (.A(_09971_),
    .B1(_09732_),
    .B2(_09749_),
    .ZN(_09972_));
 AOI21_X1 _28838_ (.A(_09972_),
    .B1(_09699_),
    .B2(_09687_),
    .ZN(_09973_));
 NOR3_X1 _28839_ (.A1(_09697_),
    .A2(_09698_),
    .A3(_09733_),
    .ZN(_09974_));
 AOI21_X1 _28840_ (.A(_09974_),
    .B1(_09820_),
    .B2(_09697_),
    .ZN(_09975_));
 OAI221_X2 _28841_ (.A(_09817_),
    .B1(_09970_),
    .B2(_09973_),
    .C1(_09975_),
    .C2(_09808_),
    .ZN(_09976_));
 NOR3_X1 _28842_ (.A1(_09811_),
    .A2(_09888_),
    .A3(_09972_),
    .ZN(_09977_));
 MUX2_X1 _28843_ (.A(net115),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(_07137_),
    .Z(_09978_));
 MUX2_X1 _28844_ (.A(_07395_),
    .B(_09978_),
    .S(_07170_),
    .Z(_09979_));
 AND2_X1 _28845_ (.A1(_09778_),
    .A2(_09979_),
    .ZN(_09980_));
 OAI21_X1 _28846_ (.A(_09887_),
    .B1(_09977_),
    .B2(_09980_),
    .ZN(_09981_));
 NOR2_X1 _28847_ (.A1(_09807_),
    .A2(_09915_),
    .ZN(_09982_));
 NAND3_X1 _28848_ (.A1(_09733_),
    .A2(_09757_),
    .A3(_09982_),
    .ZN(_09983_));
 NOR2_X4 _28849_ (.A1(_09750_),
    .A2(_09809_),
    .ZN(_09984_));
 OAI21_X1 _28850_ (.A(_09979_),
    .B1(_09984_),
    .B2(_09950_),
    .ZN(_09985_));
 NAND4_X2 _28851_ (.A1(_09976_),
    .A2(_09981_),
    .A3(_09983_),
    .A4(_09985_),
    .ZN(_09986_));
 MUX2_X1 _28852_ (.A(_12034_),
    .B(_09986_),
    .S(_09865_),
    .Z(_01549_));
 NAND2_X1 _28853_ (.A1(_09681_),
    .A2(_09820_),
    .ZN(_09987_));
 NAND3_X1 _28854_ (.A1(_09775_),
    .A2(_09860_),
    .A3(_09987_),
    .ZN(_09988_));
 MUX2_X1 _28855_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(_03978_),
    .Z(_09989_));
 MUX2_X2 _28856_ (.A(_07400_),
    .B(_09989_),
    .S(_07169_),
    .Z(_09990_));
 AOI21_X1 _28857_ (.A(_09686_),
    .B1(_09820_),
    .B2(_09990_),
    .ZN(_09991_));
 NOR2_X1 _28858_ (.A1(_09691_),
    .A2(_09991_),
    .ZN(_09992_));
 AOI21_X1 _28859_ (.A(_09992_),
    .B1(_09860_),
    .B2(_09719_),
    .ZN(_09993_));
 OAI21_X1 _28860_ (.A(_09988_),
    .B1(_09993_),
    .B2(_09772_),
    .ZN(_09994_));
 OAI21_X1 _28861_ (.A(_09816_),
    .B1(_09970_),
    .B2(_09994_),
    .ZN(_09995_));
 AOI21_X1 _28862_ (.A(_09693_),
    .B1(_09995_),
    .B2(_09695_),
    .ZN(_09996_));
 NOR2_X1 _28863_ (.A1(_09860_),
    .A2(_09996_),
    .ZN(_09997_));
 OAI21_X1 _28864_ (.A(_09752_),
    .B1(_09990_),
    .B2(_09695_),
    .ZN(_09998_));
 AOI21_X1 _28865_ (.A(_09997_),
    .B1(_09998_),
    .B2(_09995_),
    .ZN(_09999_));
 NAND2_X1 _28866_ (.A1(_09777_),
    .A2(_09990_),
    .ZN(_10000_));
 AOI22_X1 _28867_ (.A1(_09811_),
    .A2(_09722_),
    .B1(_09860_),
    .B2(_09842_),
    .ZN(_10001_));
 OAI21_X1 _28868_ (.A(_10000_),
    .B1(_10001_),
    .B2(_09808_),
    .ZN(_10002_));
 AOI22_X1 _28869_ (.A1(_09798_),
    .A2(_09999_),
    .B1(_10002_),
    .B2(_09887_),
    .ZN(_10003_));
 AOI21_X1 _28870_ (.A(_09999_),
    .B1(_09990_),
    .B2(_09798_),
    .ZN(_10004_));
 OAI21_X1 _28871_ (.A(_10003_),
    .B1(_10004_),
    .B2(_09800_),
    .ZN(_10005_));
 MUX2_X1 _28872_ (.A(_11989_),
    .B(_10005_),
    .S(_09865_),
    .Z(_01550_));
 NAND2_X2 _28873_ (.A1(_09772_),
    .A2(_09775_),
    .ZN(_10006_));
 AOI21_X1 _28874_ (.A(_09766_),
    .B1(_10006_),
    .B2(_09687_),
    .ZN(_10007_));
 OAI21_X1 _28875_ (.A(_09726_),
    .B1(_09982_),
    .B2(_10007_),
    .ZN(_10008_));
 INV_X1 _28876_ (.A(_09726_),
    .ZN(_10009_));
 MUX2_X1 _28877_ (.A(_10009_),
    .B(_09762_),
    .S(_09698_),
    .Z(_10010_));
 AOI21_X1 _28878_ (.A(_09769_),
    .B1(_09771_),
    .B2(_10010_),
    .ZN(_10011_));
 MUX2_X1 _28879_ (.A(net117),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(_07137_),
    .Z(_10012_));
 MUX2_X1 _28880_ (.A(_07402_),
    .B(_10012_),
    .S(_07170_),
    .Z(_10013_));
 AOI21_X1 _28881_ (.A(_10011_),
    .B1(_10013_),
    .B2(_09984_),
    .ZN(_10014_));
 NOR2_X1 _28882_ (.A1(_09891_),
    .A2(_10013_),
    .ZN(_10015_));
 OAI21_X1 _28883_ (.A(_09861_),
    .B1(_10013_),
    .B2(_09676_),
    .ZN(_10016_));
 OAI21_X1 _28884_ (.A(_10016_),
    .B1(_09861_),
    .B2(_10009_),
    .ZN(_10017_));
 AOI21_X1 _28885_ (.A(_09970_),
    .B1(_10017_),
    .B2(_09818_),
    .ZN(_10018_));
 OAI221_X2 _28886_ (.A(_10008_),
    .B1(_10014_),
    .B2(_10015_),
    .C1(_10018_),
    .C2(_09832_),
    .ZN(_10019_));
 MUX2_X1 _28887_ (.A(_12041_),
    .B(_10019_),
    .S(_09865_),
    .Z(_01551_));
 MUX2_X1 _28888_ (.A(net118),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(_07137_),
    .Z(_10020_));
 MUX2_X2 _28889_ (.A(_07404_),
    .B(_10020_),
    .S(_07170_),
    .Z(_10021_));
 OAI21_X1 _28890_ (.A(_09752_),
    .B1(_10021_),
    .B2(_09695_),
    .ZN(_10022_));
 OAI21_X1 _28891_ (.A(_09719_),
    .B1(_09775_),
    .B2(_09722_),
    .ZN(_10023_));
 NAND3_X1 _28892_ (.A1(_09775_),
    .A2(_09722_),
    .A3(_09819_),
    .ZN(_10024_));
 AOI21_X1 _28893_ (.A(_09772_),
    .B1(_10023_),
    .B2(_10024_),
    .ZN(_10025_));
 NAND2_X2 _28894_ (.A1(_09755_),
    .A2(_09839_),
    .ZN(_10026_));
 OAI21_X1 _28895_ (.A(_10026_),
    .B1(_09839_),
    .B2(_09853_),
    .ZN(_10027_));
 AOI221_X2 _28896_ (.A(_10025_),
    .B1(_10027_),
    .B2(_09838_),
    .C1(_09763_),
    .C2(_09848_),
    .ZN(_10028_));
 OAI21_X1 _28897_ (.A(_10022_),
    .B1(_10028_),
    .B2(_09766_),
    .ZN(_10029_));
 OAI21_X1 _28898_ (.A(_10029_),
    .B1(_09722_),
    .B2(_09808_),
    .ZN(_10030_));
 AOI22_X2 _28899_ (.A1(_09771_),
    .A2(_09763_),
    .B1(_10021_),
    .B2(_09778_),
    .ZN(_10031_));
 OAI21_X1 _28900_ (.A(_10021_),
    .B1(_09821_),
    .B2(_09798_),
    .ZN(_10032_));
 OAI221_X2 _28901_ (.A(_10030_),
    .B1(_10031_),
    .B2(_09769_),
    .C1(_09800_),
    .C2(_10032_),
    .ZN(_10033_));
 MUX2_X1 _28902_ (.A(_11992_),
    .B(_10033_),
    .S(_09865_),
    .Z(_01552_));
 NAND2_X4 _28903_ (.A1(_09694_),
    .A2(_09817_),
    .ZN(_10034_));
 NAND2_X1 _28904_ (.A1(_09807_),
    .A2(_09841_),
    .ZN(_10035_));
 AOI21_X1 _28905_ (.A(_10035_),
    .B1(_09839_),
    .B2(_09699_),
    .ZN(_10036_));
 OAI21_X1 _28906_ (.A(_09771_),
    .B1(_09775_),
    .B2(_09755_),
    .ZN(_10037_));
 INV_X1 _28907_ (.A(_10037_),
    .ZN(_10038_));
 NAND2_X2 _28908_ (.A1(_09755_),
    .A2(_09851_),
    .ZN(_10039_));
 NAND2_X1 _28909_ (.A1(_07137_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .ZN(_10040_));
 NAND2_X1 _28910_ (.A1(_09749_),
    .A2(net119),
    .ZN(_10041_));
 AOI21_X1 _28911_ (.A(_03981_),
    .B1(_10040_),
    .B2(_10041_),
    .ZN(_10042_));
 AOI21_X2 _28912_ (.A(_10042_),
    .B1(_07405_),
    .B2(_03981_),
    .ZN(_10043_));
 AOI21_X1 _28913_ (.A(_10039_),
    .B1(_10043_),
    .B2(_09805_),
    .ZN(_10044_));
 INV_X1 _28914_ (.A(_10026_),
    .ZN(_10045_));
 AOI22_X1 _28915_ (.A1(_09697_),
    .A2(_09841_),
    .B1(_09872_),
    .B2(_10045_),
    .ZN(_10046_));
 NOR2_X1 _28916_ (.A1(_09823_),
    .A2(_10046_),
    .ZN(_10047_));
 NOR4_X2 _28917_ (.A1(_10036_),
    .A2(_10038_),
    .A3(_10044_),
    .A4(_10047_),
    .ZN(_10048_));
 AOI21_X4 _28918_ (.A(_09984_),
    .B1(_09777_),
    .B2(_09884_),
    .ZN(_10049_));
 AOI22_X2 _28919_ (.A1(_09884_),
    .A2(_09891_),
    .B1(_09752_),
    .B2(_09776_),
    .ZN(_10050_));
 OAI222_X2 _28920_ (.A1(_10034_),
    .A2(_10048_),
    .B1(_10049_),
    .B2(_10043_),
    .C1(_10050_),
    .C2(_09676_),
    .ZN(_10051_));
 MUX2_X1 _28921_ (.A(_10873_),
    .B(_10051_),
    .S(_09865_),
    .Z(_01553_));
 MUX2_X1 _28922_ (.A(_09841_),
    .B(_09710_),
    .S(_09697_),
    .Z(_10052_));
 NAND3_X1 _28923_ (.A1(_09776_),
    .A2(_09752_),
    .A3(_10052_),
    .ZN(_10053_));
 AOI221_X2 _28924_ (.A(_09769_),
    .B1(_09776_),
    .B2(_10009_),
    .C1(_09867_),
    .C2(_09693_),
    .ZN(_10054_));
 NOR2_X1 _28925_ (.A1(_09984_),
    .A2(_10054_),
    .ZN(_10055_));
 MUX2_X1 _28926_ (.A(net120),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(_07136_),
    .Z(_10056_));
 MUX2_X1 _28927_ (.A(_07335_),
    .B(_10056_),
    .S(_07170_),
    .Z(_10057_));
 AOI21_X1 _28928_ (.A(_10057_),
    .B1(_10054_),
    .B2(_09891_),
    .ZN(_10058_));
 NAND3_X1 _28929_ (.A1(_09807_),
    .A2(_09823_),
    .A3(_09710_),
    .ZN(_10059_));
 AOI21_X1 _28930_ (.A(_10038_),
    .B1(_09842_),
    .B2(_09726_),
    .ZN(_10060_));
 INV_X1 _28931_ (.A(_10039_),
    .ZN(_10061_));
 OAI21_X1 _28932_ (.A(_10061_),
    .B1(_10057_),
    .B2(_09762_),
    .ZN(_10062_));
 NAND3_X1 _28933_ (.A1(_10059_),
    .A2(_10060_),
    .A3(_10062_),
    .ZN(_10063_));
 OAI21_X1 _28934_ (.A(_10026_),
    .B1(_09839_),
    .B2(_10009_),
    .ZN(_10064_));
 AOI21_X1 _28935_ (.A(_10063_),
    .B1(_10064_),
    .B2(_09838_),
    .ZN(_10065_));
 OAI221_X2 _28936_ (.A(_10053_),
    .B1(_10055_),
    .B2(_10058_),
    .C1(_10034_),
    .C2(_10065_),
    .ZN(_10066_));
 BUF_X4 _28937_ (.A(_07180_),
    .Z(_10067_));
 MUX2_X1 _28938_ (.A(_10874_),
    .B(_10066_),
    .S(_10067_),
    .Z(_01554_));
 MUX2_X1 _28939_ (.A(net121),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(_07136_),
    .Z(_10068_));
 MUX2_X2 _28940_ (.A(_07336_),
    .B(_10068_),
    .S(_07169_),
    .Z(_10069_));
 NOR2_X1 _28941_ (.A1(_09762_),
    .A2(_10069_),
    .ZN(_10070_));
 NOR2_X1 _28942_ (.A1(_09842_),
    .A2(_09848_),
    .ZN(_10071_));
 OAI221_X1 _28943_ (.A(_10037_),
    .B1(_10039_),
    .B2(_10070_),
    .C1(_10071_),
    .C2(_09853_),
    .ZN(_10072_));
 OAI21_X1 _28944_ (.A(_10026_),
    .B1(_09839_),
    .B2(_09972_),
    .ZN(_10073_));
 AOI21_X1 _28945_ (.A(_10072_),
    .B1(_10073_),
    .B2(_09838_),
    .ZN(_10074_));
 NOR2_X1 _28946_ (.A1(_10034_),
    .A2(_10074_),
    .ZN(_10075_));
 AOI21_X1 _28947_ (.A(_09800_),
    .B1(_09797_),
    .B2(_10069_),
    .ZN(_10076_));
 MUX2_X1 _28948_ (.A(_09704_),
    .B(_09972_),
    .S(_09719_),
    .Z(_10077_));
 OAI21_X1 _28949_ (.A(_09809_),
    .B1(_10077_),
    .B2(_09823_),
    .ZN(_10078_));
 OAI21_X1 _28950_ (.A(_10078_),
    .B1(_10069_),
    .B2(_09695_),
    .ZN(_10079_));
 AOI21_X1 _28951_ (.A(_10076_),
    .B1(_10079_),
    .B2(_09798_),
    .ZN(_10080_));
 NOR2_X1 _28952_ (.A1(_10075_),
    .A2(_10080_),
    .ZN(_10081_));
 AOI22_X1 _28953_ (.A1(_09703_),
    .A2(_09693_),
    .B1(_10069_),
    .B2(_09778_),
    .ZN(_10082_));
 AOI21_X1 _28954_ (.A(_10081_),
    .B1(_10082_),
    .B2(_09887_),
    .ZN(_10083_));
 MUX2_X1 _28955_ (.A(_10500_),
    .B(_10083_),
    .S(_10067_),
    .Z(_01555_));
 MUX2_X1 _28956_ (.A(net122),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(_07136_),
    .Z(_10084_));
 MUX2_X1 _28957_ (.A(_07337_),
    .B(_10084_),
    .S(_07169_),
    .Z(_10085_));
 NAND2_X1 _28958_ (.A1(_09984_),
    .A2(_10085_),
    .ZN(_10086_));
 AOI22_X2 _28959_ (.A1(_09707_),
    .A2(_09693_),
    .B1(_10085_),
    .B2(_09778_),
    .ZN(_10087_));
 OAI21_X1 _28960_ (.A(_09757_),
    .B1(_09707_),
    .B2(_09691_),
    .ZN(_10088_));
 AOI221_X2 _28961_ (.A(_09818_),
    .B1(_10088_),
    .B2(_09772_),
    .C1(_09691_),
    .C2(_09676_),
    .ZN(_10089_));
 OR2_X1 _28962_ (.A1(_09762_),
    .A2(_10085_),
    .ZN(_10090_));
 INV_X1 _28963_ (.A(_09860_),
    .ZN(_10091_));
 OAI21_X1 _28964_ (.A(_10026_),
    .B1(_09839_),
    .B2(_10091_),
    .ZN(_10092_));
 AOI221_X2 _28965_ (.A(_10089_),
    .B1(_10090_),
    .B2(_10061_),
    .C1(_10092_),
    .C2(_09838_),
    .ZN(_10093_));
 OAI221_X2 _28966_ (.A(_10086_),
    .B1(_10087_),
    .B2(_09769_),
    .C1(_10034_),
    .C2(_10093_),
    .ZN(_10094_));
 MUX2_X1 _28967_ (.A(net305),
    .B(_10094_),
    .S(_10067_),
    .Z(_01556_));
 NAND2_X1 _28968_ (.A1(_10502_),
    .A2(_07253_),
    .ZN(_10095_));
 MUX2_X1 _28969_ (.A(net123),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(_07136_),
    .Z(_10096_));
 MUX2_X2 _28970_ (.A(_07338_),
    .B(_10096_),
    .S(_07170_),
    .Z(_10097_));
 AOI22_X1 _28971_ (.A1(_09805_),
    .A2(_09693_),
    .B1(_10097_),
    .B2(_09777_),
    .ZN(_10098_));
 NOR2_X1 _28972_ (.A1(_09769_),
    .A2(_10098_),
    .ZN(_10099_));
 OAI21_X1 _28973_ (.A(_09756_),
    .B1(_09698_),
    .B2(_09771_),
    .ZN(_10100_));
 NOR2_X1 _28974_ (.A1(_09762_),
    .A2(_10097_),
    .ZN(_10101_));
 OAI221_X2 _28975_ (.A(_10100_),
    .B1(_10101_),
    .B2(_10039_),
    .C1(_10006_),
    .C2(_09762_),
    .ZN(_10102_));
 AOI221_X2 _28976_ (.A(_10099_),
    .B1(_10097_),
    .B2(_09984_),
    .C1(_09817_),
    .C2(_10102_),
    .ZN(_10103_));
 OAI21_X1 _28977_ (.A(_10095_),
    .B1(_10103_),
    .B2(_09783_),
    .ZN(_01557_));
 INV_X1 _28978_ (.A(_09718_),
    .ZN(_10104_));
 AOI21_X1 _28979_ (.A(_09738_),
    .B1(_09756_),
    .B2(_10104_),
    .ZN(_10105_));
 NAND3_X1 _28980_ (.A1(_09818_),
    .A2(_09752_),
    .A3(_10105_),
    .ZN(_10106_));
 OR2_X1 _28981_ (.A1(_09868_),
    .A2(_09832_),
    .ZN(_10107_));
 AND2_X1 _28982_ (.A1(_10049_),
    .A2(_10107_),
    .ZN(_10108_));
 OAI221_X2 _28983_ (.A(_10106_),
    .B1(_09908_),
    .B2(_09832_),
    .C1(_09965_),
    .C2(_10108_),
    .ZN(_10109_));
 MUX2_X1 _28984_ (.A(\id_stage_i.controller_i.instr_i[2] ),
    .B(_10109_),
    .S(_10067_),
    .Z(_01558_));
 NAND2_X1 _28985_ (.A1(_07136_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .ZN(_10110_));
 NAND2_X1 _28986_ (.A1(_09749_),
    .A2(net125),
    .ZN(_10111_));
 AOI21_X2 _28987_ (.A(_03963_),
    .B1(_10110_),
    .B2(_10111_),
    .ZN(_10112_));
 AOI21_X4 _28988_ (.A(_10112_),
    .B1(_07339_),
    .B2(_03981_),
    .ZN(_10113_));
 NAND2_X1 _28989_ (.A1(_09820_),
    .A2(_10113_),
    .ZN(_10114_));
 AOI21_X1 _28990_ (.A(_09762_),
    .B1(_09763_),
    .B2(_09779_),
    .ZN(_10115_));
 OAI221_X2 _28991_ (.A(_10114_),
    .B1(_10115_),
    .B2(_09755_),
    .C1(_09763_),
    .C2(_09805_),
    .ZN(_10116_));
 AOI221_X2 _28992_ (.A(_09698_),
    .B1(_09835_),
    .B2(_10116_),
    .C1(_09704_),
    .C2(_09807_),
    .ZN(_10117_));
 AOI21_X2 _28993_ (.A(_10117_),
    .B1(_09756_),
    .B2(_09699_),
    .ZN(_10118_));
 OAI22_X4 _28994_ (.A1(_10049_),
    .A2(_10113_),
    .B1(_10118_),
    .B2(_10034_),
    .ZN(_10119_));
 MUX2_X1 _28995_ (.A(_10498_),
    .B(_10119_),
    .S(_10067_),
    .Z(_01559_));
 NAND2_X1 _28996_ (.A1(_07137_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .ZN(_10120_));
 NAND2_X1 _28997_ (.A1(_09749_),
    .A2(net126),
    .ZN(_10121_));
 AOI21_X1 _28998_ (.A(_03981_),
    .B1(_10120_),
    .B2(_10121_),
    .ZN(_10122_));
 AOI21_X2 _28999_ (.A(_10122_),
    .B1(_07340_),
    .B2(_03981_),
    .ZN(_10123_));
 AOI21_X1 _29000_ (.A(_10039_),
    .B1(_10123_),
    .B2(_09805_),
    .ZN(_10124_));
 AOI21_X1 _29001_ (.A(_10124_),
    .B1(_09760_),
    .B2(_09756_),
    .ZN(_10125_));
 OAI22_X2 _29002_ (.A1(_10049_),
    .A2(_10123_),
    .B1(_10125_),
    .B2(_10034_),
    .ZN(_10126_));
 MUX2_X1 _29003_ (.A(_10509_),
    .B(_10126_),
    .S(_10067_),
    .Z(_01560_));
 OAI22_X1 _29004_ (.A1(_09766_),
    .A2(_10006_),
    .B1(_10108_),
    .B2(_09972_),
    .ZN(_10127_));
 MUX2_X1 _29005_ (.A(_10341_),
    .B(_10127_),
    .S(_10067_),
    .Z(_01561_));
 AOI21_X1 _29006_ (.A(_09807_),
    .B1(_09697_),
    .B2(_09828_),
    .ZN(_10128_));
 AOI21_X1 _29007_ (.A(_09699_),
    .B1(_09885_),
    .B2(_10105_),
    .ZN(_10129_));
 OAI221_X1 _29008_ (.A(_09800_),
    .B1(_09860_),
    .B2(_10128_),
    .C1(_10129_),
    .C2(_09808_),
    .ZN(_10130_));
 AOI21_X1 _29009_ (.A(_09797_),
    .B1(_09697_),
    .B2(_09820_),
    .ZN(_10131_));
 OAI221_X1 _29010_ (.A(_09795_),
    .B1(_09798_),
    .B2(_10071_),
    .C1(_10131_),
    .C2(_09860_),
    .ZN(_10132_));
 AND3_X1 _29011_ (.A1(_07180_),
    .A2(_10130_),
    .A3(_10132_),
    .ZN(_10133_));
 AOI21_X1 _29012_ (.A(_10133_),
    .B1(_09783_),
    .B2(_10372_),
    .ZN(_01562_));
 OAI21_X1 _29013_ (.A(_09861_),
    .B1(_09676_),
    .B2(_09726_),
    .ZN(_10134_));
 AOI21_X1 _29014_ (.A(_09811_),
    .B1(_09823_),
    .B2(_10134_),
    .ZN(_10135_));
 OAI221_X1 _29015_ (.A(_09817_),
    .B1(_09757_),
    .B2(_09839_),
    .C1(_10135_),
    .C2(_09808_),
    .ZN(_10136_));
 AOI21_X1 _29016_ (.A(_09800_),
    .B1(_09797_),
    .B2(_09726_),
    .ZN(_10137_));
 NOR2_X1 _29017_ (.A1(_09826_),
    .A2(_10137_),
    .ZN(_10138_));
 AOI21_X1 _29018_ (.A(_09808_),
    .B1(_09823_),
    .B2(_09828_),
    .ZN(_10139_));
 OAI21_X1 _29019_ (.A(_10138_),
    .B1(_10139_),
    .B2(_09726_),
    .ZN(_10140_));
 AND3_X1 _29020_ (.A1(_07180_),
    .A2(_10136_),
    .A3(_10140_),
    .ZN(_10141_));
 AOI21_X1 _29021_ (.A(_10141_),
    .B1(_09783_),
    .B2(_10289_),
    .ZN(_01563_));
 NAND2_X1 _29022_ (.A1(_09750_),
    .A2(_09698_),
    .ZN(_10142_));
 NOR2_X1 _29023_ (.A1(_09800_),
    .A2(_10142_),
    .ZN(_10143_));
 AOI21_X1 _29024_ (.A(_10143_),
    .B1(_09982_),
    .B2(_09739_),
    .ZN(_10144_));
 OAI222_X2 _29025_ (.A1(_09766_),
    .A2(_10006_),
    .B1(_10108_),
    .B2(_09853_),
    .C1(_09811_),
    .C2(_10144_),
    .ZN(_10145_));
 MUX2_X1 _29026_ (.A(_10299_),
    .B(_10145_),
    .S(_10067_),
    .Z(_01564_));
 NOR2_X1 _29027_ (.A1(_10104_),
    .A2(_09957_),
    .ZN(_10146_));
 OAI21_X1 _29028_ (.A(_09800_),
    .B1(_09828_),
    .B2(_10146_),
    .ZN(_10147_));
 AOI21_X1 _29029_ (.A(_09872_),
    .B1(_09835_),
    .B2(_09710_),
    .ZN(_10148_));
 NOR2_X1 _29030_ (.A1(_09698_),
    .A2(_10148_),
    .ZN(_10149_));
 AOI21_X1 _29031_ (.A(_10149_),
    .B1(_09842_),
    .B2(_09756_),
    .ZN(_10150_));
 OAI21_X1 _29032_ (.A(_10147_),
    .B1(_10150_),
    .B2(_09798_),
    .ZN(_10151_));
 OAI21_X1 _29033_ (.A(_09835_),
    .B1(_09956_),
    .B2(_09698_),
    .ZN(_10152_));
 AOI21_X1 _29034_ (.A(_09745_),
    .B1(_09797_),
    .B2(_10152_),
    .ZN(_10153_));
 AOI21_X1 _29035_ (.A(_09797_),
    .B1(_09719_),
    .B2(_10006_),
    .ZN(_10154_));
 NOR2_X1 _29036_ (.A1(_10153_),
    .A2(_10154_),
    .ZN(_10155_));
 OAI21_X1 _29037_ (.A(_09884_),
    .B1(_09687_),
    .B2(_09965_),
    .ZN(_10156_));
 OAI22_X1 _29038_ (.A1(_10151_),
    .A2(_10155_),
    .B1(_10156_),
    .B2(_09778_),
    .ZN(_10157_));
 AOI21_X1 _29039_ (.A(_09710_),
    .B1(_10151_),
    .B2(_10156_),
    .ZN(_10158_));
 NOR2_X1 _29040_ (.A1(_10157_),
    .A2(_10158_),
    .ZN(_10159_));
 MUX2_X1 _29041_ (.A(_10902_),
    .B(_10159_),
    .S(_10067_),
    .Z(_01565_));
 NAND3_X1 _29042_ (.A1(_09817_),
    .A2(_09733_),
    .A3(_09842_),
    .ZN(_10160_));
 AOI21_X1 _29043_ (.A(_10155_),
    .B1(_09818_),
    .B2(_09817_),
    .ZN(_10161_));
 AOI22_X1 _29044_ (.A1(_09778_),
    .A2(_09703_),
    .B1(_09733_),
    .B2(_09771_),
    .ZN(_10162_));
 OAI221_X1 _29045_ (.A(_10160_),
    .B1(_10161_),
    .B2(_09704_),
    .C1(_10162_),
    .C2(_09769_),
    .ZN(_10163_));
 MUX2_X1 _29046_ (.A(_10394_),
    .B(_10163_),
    .S(_10067_),
    .Z(_01566_));
 NAND2_X1 _29047_ (.A1(_06224_),
    .A2(_07253_),
    .ZN(_10164_));
 INV_X1 _29048_ (.A(_09707_),
    .ZN(_10165_));
 AOI22_X1 _29049_ (.A1(_09811_),
    .A2(_09860_),
    .B1(_09842_),
    .B2(_09722_),
    .ZN(_10166_));
 OAI221_X1 _29050_ (.A(_09887_),
    .B1(_09891_),
    .B2(_10165_),
    .C1(_10166_),
    .C2(_09808_),
    .ZN(_10167_));
 AOI21_X1 _29051_ (.A(_09798_),
    .B1(_10006_),
    .B2(_09795_),
    .ZN(_10168_));
 AOI21_X1 _29052_ (.A(_09811_),
    .B1(_09810_),
    .B2(_10142_),
    .ZN(_10169_));
 OAI33_X1 _29053_ (.A1(_09811_),
    .A2(_10091_),
    .A3(_10142_),
    .B1(_10168_),
    .B2(_10169_),
    .B3(_10165_),
    .ZN(_10170_));
 OAI21_X1 _29054_ (.A(_10167_),
    .B1(_10170_),
    .B2(_09887_),
    .ZN(_10171_));
 OAI21_X1 _29055_ (.A(_10164_),
    .B1(_10171_),
    .B2(_09783_),
    .ZN(_01567_));
 CLKBUF_X3 _29056_ (.A(_07180_),
    .Z(_10172_));
 MUX2_X1 _29057_ (.A(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .B(_09795_),
    .S(_10172_),
    .Z(_01568_));
 MUX2_X1 _29058_ (.A(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .B(_09805_),
    .S(_10172_),
    .Z(_01569_));
 MUX2_X1 _29059_ (.A(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .B(_09763_),
    .S(_10172_),
    .Z(_01570_));
 MUX2_X1 _29060_ (.A(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .B(_09756_),
    .S(_10172_),
    .Z(_01571_));
 MUX2_X1 _29061_ (.A(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .B(_09808_),
    .S(_10172_),
    .Z(_01572_));
 MUX2_X1 _29062_ (.A(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .B(_09699_),
    .S(_10172_),
    .Z(_01573_));
 MUX2_X1 _29063_ (.A(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .B(_09697_),
    .S(_10172_),
    .Z(_01574_));
 MUX2_X1 _29064_ (.A(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .B(_09798_),
    .S(_10172_),
    .Z(_01575_));
 MUX2_X1 _29065_ (.A(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .B(_09841_),
    .S(_10172_),
    .Z(_01576_));
 MUX2_X1 _29066_ (.A(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .B(_09733_),
    .S(_10172_),
    .Z(_01577_));
 BUF_X4 _29067_ (.A(_07180_),
    .Z(_10173_));
 MUX2_X1 _29068_ (.A(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .B(_09860_),
    .S(_10173_),
    .Z(_01578_));
 MUX2_X1 _29069_ (.A(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .B(_09726_),
    .S(_10173_),
    .Z(_01579_));
 MUX2_X1 _29070_ (.A(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .B(_09722_),
    .S(_10173_),
    .Z(_01580_));
 MUX2_X1 _29071_ (.A(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .B(_09710_),
    .S(_10173_),
    .Z(_01581_));
 MUX2_X1 _29072_ (.A(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .B(_09703_),
    .S(_10173_),
    .Z(_01582_));
 MUX2_X1 _29073_ (.A(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .B(_09707_),
    .S(_10173_),
    .Z(_01583_));
 MUX2_X1 _29074_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(\cs_registers_i.pc_if_i[10] ),
    .S(_10173_),
    .Z(_01584_));
 MUX2_X1 _29075_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_07178_),
    .S(_10173_),
    .Z(_01585_));
 MUX2_X1 _29076_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(_07199_),
    .S(_10173_),
    .Z(_01586_));
 MUX2_X1 _29077_ (.A(_12076_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .S(_10173_),
    .Z(_01587_));
 CLKBUF_X3 _29078_ (.A(_07180_),
    .Z(_10174_));
 MUX2_X1 _29079_ (.A(_12179_),
    .B(\cs_registers_i.pc_if_i[14] ),
    .S(_10174_),
    .Z(_01588_));
 MUX2_X1 _29080_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_07222_),
    .S(_10174_),
    .Z(_01589_));
 MUX2_X1 _29081_ (.A(\cs_registers_i.pc_id_i[16] ),
    .B(\cs_registers_i.pc_if_i[16] ),
    .S(_10174_),
    .Z(_01590_));
 MUX2_X1 _29082_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(\cs_registers_i.pc_if_i[17] ),
    .S(_10174_),
    .Z(_01591_));
 MUX2_X1 _29083_ (.A(\cs_registers_i.pc_id_i[18] ),
    .B(_07235_),
    .S(_10174_),
    .Z(_01592_));
 MUX2_X1 _29084_ (.A(_12590_),
    .B(_07241_),
    .S(_10174_),
    .Z(_01593_));
 MUX2_X1 _29085_ (.A(_03981_),
    .B(_10675_),
    .S(_07253_),
    .Z(_01594_));
 MUX2_X1 _29086_ (.A(_12685_),
    .B(_07249_),
    .S(_10174_),
    .Z(_01595_));
 MUX2_X1 _29087_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(\cs_registers_i.pc_if_i[21] ),
    .S(_10174_),
    .Z(_01596_));
 MUX2_X1 _29088_ (.A(\cs_registers_i.pc_id_i[22] ),
    .B(_07259_),
    .S(_10174_),
    .Z(_01597_));
 MUX2_X1 _29089_ (.A(_12935_),
    .B(_07263_),
    .S(_10174_),
    .Z(_01598_));
 CLKBUF_X3 _29090_ (.A(_07179_),
    .Z(_10175_));
 MUX2_X1 _29091_ (.A(_13024_),
    .B(\cs_registers_i.pc_if_i[24] ),
    .S(_10175_),
    .Z(_01599_));
 MUX2_X1 _29092_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(\cs_registers_i.pc_if_i[25] ),
    .S(_10175_),
    .Z(_01600_));
 MUX2_X1 _29093_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(_07281_),
    .S(_10175_),
    .Z(_01601_));
 MUX2_X1 _29094_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(_07285_),
    .S(_10175_),
    .Z(_01602_));
 MUX2_X1 _29095_ (.A(\cs_registers_i.pc_id_i[28] ),
    .B(\cs_registers_i.pc_if_i[28] ),
    .S(_10175_),
    .Z(_01603_));
 MUX2_X1 _29096_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(\cs_registers_i.pc_if_i[29] ),
    .S(_10175_),
    .Z(_01604_));
 MUX2_X1 _29097_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(\cs_registers_i.pc_if_i[2] ),
    .S(_10175_),
    .Z(_01605_));
 MUX2_X1 _29098_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(\cs_registers_i.pc_if_i[30] ),
    .S(_10175_),
    .Z(_01606_));
 MUX2_X1 _29099_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(\cs_registers_i.pc_if_i[31] ),
    .S(_10175_),
    .Z(_01607_));
 MUX2_X1 _29100_ (.A(_11517_),
    .B(_07181_),
    .S(_10175_),
    .Z(_01608_));
 MUX2_X1 _29101_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(_07186_),
    .S(_07193_),
    .Z(_01609_));
 MUX2_X1 _29102_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_07187_),
    .S(_07193_),
    .Z(_01610_));
 MUX2_X1 _29103_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(\cs_registers_i.pc_if_i[6] ),
    .S(_07193_),
    .Z(_01611_));
 MUX2_X1 _29104_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_07185_),
    .S(_07193_),
    .Z(_01612_));
 MUX2_X1 _29105_ (.A(_11788_),
    .B(\cs_registers_i.pc_if_i[8] ),
    .S(_07193_),
    .Z(_01613_));
 MUX2_X1 _29106_ (.A(_11826_),
    .B(_07184_),
    .S(_07193_),
    .Z(_01614_));
 NAND2_X2 _29107_ (.A1(_00133_),
    .A2(_04162_),
    .ZN(net254));
 NOR4_X1 _29108_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_04155_),
    .A3(_07425_),
    .A4(_06287_),
    .ZN(_10176_));
 OAI21_X1 _29109_ (.A(_10176_),
    .B1(_06286_),
    .B2(_03436_),
    .ZN(_10177_));
 OR2_X1 _29110_ (.A1(net254),
    .A2(_10177_),
    .ZN(core_busy_d));
 AND2_X1 _29111_ (.A1(clknet_1_0__leaf_clk_i),
    .A2(\core_clock_gate_i.en_latch ),
    .ZN(clk));
 NOR2_X1 _29112_ (.A1(_10477_),
    .A2(_03619_),
    .ZN(_10178_));
 AOI21_X1 _29113_ (.A(_10178_),
    .B1(_16086_),
    .B2(_10477_),
    .ZN(_10179_));
 MUX2_X2 _29114_ (.A(_16087_),
    .B(_10179_),
    .S(_07447_),
    .Z(net186));
 MUX2_X1 _29115_ (.A(_16101_),
    .B(_16091_),
    .S(_10477_),
    .Z(_10180_));
 MUX2_X2 _29116_ (.A(_16089_),
    .B(_10180_),
    .S(_07447_),
    .Z(net187));
 NAND2_X1 _29117_ (.A1(_16097_),
    .A2(_07475_),
    .ZN(_10181_));
 INV_X1 _29118_ (.A(_07446_),
    .ZN(_10182_));
 OAI21_X1 _29119_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B1(_07447_),
    .B2(_10182_),
    .ZN(_10183_));
 NAND3_X1 _29120_ (.A1(_10477_),
    .A2(_16094_),
    .A3(_07447_),
    .ZN(_10184_));
 OAI21_X1 _29121_ (.A(_10184_),
    .B1(_07447_),
    .B2(_16093_),
    .ZN(_10185_));
 OAI21_X1 _29122_ (.A(_10183_),
    .B1(_10185_),
    .B2(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_10186_));
 NAND2_X2 _29123_ (.A1(_10181_),
    .A2(_10186_),
    .ZN(net188));
 MUX2_X1 _29124_ (.A(_07446_),
    .B(_16088_),
    .S(_10477_),
    .Z(_10187_));
 MUX2_X2 _29125_ (.A(_16085_),
    .B(_10187_),
    .S(_07447_),
    .Z(net189));
 BUF_X2 _29126_ (.A(_16099_),
    .Z(_10188_));
 BUF_X4 _29127_ (.A(_10188_),
    .Z(_10189_));
 BUF_X2 _29128_ (.A(_16103_),
    .Z(_10190_));
 AOI22_X1 _29129_ (.A1(_10189_),
    .A2(_12316_),
    .B1(_12985_),
    .B2(_10190_),
    .ZN(_10191_));
 OAI21_X1 _29130_ (.A(_10191_),
    .B1(_11241_),
    .B2(_10182_),
    .ZN(_10192_));
 NOR2_X1 _29131_ (.A1(_03619_),
    .A2(_10192_),
    .ZN(_10193_));
 AOI21_X4 _29132_ (.A(_10193_),
    .B1(_03660_),
    .B2(_03619_),
    .ZN(net191));
 BUF_X8 _29133_ (.A(_03620_),
    .Z(_10194_));
 NOR2_X1 _29134_ (.A1(_10194_),
    .A2(_03736_),
    .ZN(_10195_));
 BUF_X4 _29135_ (.A(_07446_),
    .Z(_10196_));
 BUF_X4 _29136_ (.A(_10196_),
    .Z(_10197_));
 BUF_X4 _29137_ (.A(_10188_),
    .Z(_10198_));
 BUF_X4 _29138_ (.A(_10190_),
    .Z(_10199_));
 AOI222_X2 _29139_ (.A1(_10197_),
    .A2(net346),
    .B1(net313),
    .B2(_10198_),
    .C1(_10199_),
    .C2(_10973_),
    .ZN(_10200_));
 AOI21_X2 _29140_ (.A(_10195_),
    .B1(_10200_),
    .B2(_16084_),
    .ZN(net192));
 NOR2_X1 _29141_ (.A1(_10194_),
    .A2(_11351_),
    .ZN(_10201_));
 AOI222_X2 _29142_ (.A1(_10197_),
    .A2(net281),
    .B1(net329),
    .B2(_10198_),
    .C1(_10199_),
    .C2(_11019_),
    .ZN(_10202_));
 AOI21_X2 _29143_ (.A(_10201_),
    .B1(_10202_),
    .B2(_16084_),
    .ZN(net193));
 CLKBUF_X3 _29144_ (.A(_03620_),
    .Z(_10203_));
 NOR2_X1 _29145_ (.A1(_10203_),
    .A2(net303),
    .ZN(_10204_));
 AOI222_X2 _29146_ (.A1(_10197_),
    .A2(net355),
    .B1(net330),
    .B2(_10198_),
    .C1(_10199_),
    .C2(_03519_),
    .ZN(_10205_));
 AOI21_X2 _29147_ (.A(_10204_),
    .B1(_10205_),
    .B2(_16084_),
    .ZN(net194));
 NOR2_X1 _29148_ (.A1(_10203_),
    .A2(_12044_),
    .ZN(_10206_));
 BUF_X4 _29149_ (.A(_10188_),
    .Z(_10207_));
 BUF_X4 _29150_ (.A(_10190_),
    .Z(_10208_));
 AOI222_X2 _29151_ (.A1(_10197_),
    .A2(net290),
    .B1(_03166_),
    .B2(_10207_),
    .C1(_10208_),
    .C2(_03696_),
    .ZN(_10209_));
 AOI21_X2 _29152_ (.A(_10206_),
    .B1(_10209_),
    .B2(_16084_),
    .ZN(net195));
 NOR2_X1 _29153_ (.A1(_10203_),
    .A2(_12144_),
    .ZN(_10210_));
 AOI222_X2 _29154_ (.A1(_10197_),
    .A2(net288),
    .B1(_03275_),
    .B2(_10207_),
    .C1(_10208_),
    .C2(_11158_),
    .ZN(_10211_));
 AOI21_X2 _29155_ (.A(_10210_),
    .B1(_10211_),
    .B2(_16084_),
    .ZN(net196));
 NOR2_X1 _29156_ (.A1(_10203_),
    .A2(net327),
    .ZN(_10212_));
 AOI222_X2 _29157_ (.A1(_10197_),
    .A2(net286),
    .B1(_03772_),
    .B2(_10207_),
    .C1(_10208_),
    .C2(_11202_),
    .ZN(_10213_));
 AOI21_X2 _29158_ (.A(_10212_),
    .B1(_10213_),
    .B2(_16084_),
    .ZN(net197));
 NAND2_X1 _29159_ (.A1(_10196_),
    .A2(_12985_),
    .ZN(_10214_));
 BUF_X4 _29160_ (.A(_10190_),
    .Z(_10215_));
 INV_X1 _29161_ (.A(_10215_),
    .ZN(_10216_));
 INV_X1 _29162_ (.A(_10189_),
    .ZN(_10217_));
 OAI221_X1 _29163_ (.A(_10214_),
    .B1(_11241_),
    .B2(_10216_),
    .C1(_10217_),
    .C2(_03660_),
    .ZN(_10218_));
 MUX2_X2 _29164_ (.A(_12316_),
    .B(_10218_),
    .S(_04153_),
    .Z(net198));
 NOR2_X1 _29165_ (.A1(_10203_),
    .A2(net344),
    .ZN(_10219_));
 AOI222_X2 _29166_ (.A1(_10198_),
    .A2(net348),
    .B1(_03727_),
    .B2(_10199_),
    .C1(net292),
    .C2(_10196_),
    .ZN(_10220_));
 AOI21_X2 _29167_ (.A(_10219_),
    .B1(_10220_),
    .B2(_16084_),
    .ZN(net199));
 NOR2_X1 _29168_ (.A1(_10203_),
    .A2(_12482_),
    .ZN(_10221_));
 AOI222_X2 _29169_ (.A1(_10198_),
    .A2(_10973_),
    .B1(_03736_),
    .B2(_10199_),
    .C1(net314),
    .C2(_10196_),
    .ZN(_10222_));
 AOI21_X2 _29170_ (.A(_10221_),
    .B1(_10222_),
    .B2(_16084_),
    .ZN(net200));
 NOR2_X1 _29171_ (.A1(_10203_),
    .A2(net281),
    .ZN(_10223_));
 AOI222_X2 _29172_ (.A1(_10198_),
    .A2(_11019_),
    .B1(_11351_),
    .B2(_10199_),
    .C1(net329),
    .C2(_10196_),
    .ZN(_10224_));
 AOI21_X2 _29173_ (.A(_10223_),
    .B1(_10224_),
    .B2(_16084_),
    .ZN(net201));
 NOR2_X1 _29174_ (.A1(_10203_),
    .A2(net348),
    .ZN(_10225_));
 AOI222_X2 _29175_ (.A1(_10197_),
    .A2(_03727_),
    .B1(net344),
    .B2(_10207_),
    .C1(net292),
    .C2(_10208_),
    .ZN(_10226_));
 BUF_X8 _29176_ (.A(_04153_),
    .Z(_10227_));
 AOI21_X2 _29177_ (.A(_10225_),
    .B1(_10226_),
    .B2(_10227_),
    .ZN(net202));
 NOR2_X1 _29178_ (.A1(_10203_),
    .A2(net355),
    .ZN(_10228_));
 AOI222_X2 _29179_ (.A1(_10198_),
    .A2(_03519_),
    .B1(net303),
    .B2(_10199_),
    .C1(net330),
    .C2(_10196_),
    .ZN(_10229_));
 AOI21_X2 _29180_ (.A(_10228_),
    .B1(_10229_),
    .B2(_10227_),
    .ZN(net203));
 NOR2_X1 _29181_ (.A1(_10203_),
    .A2(net290),
    .ZN(_10230_));
 AOI222_X2 _29182_ (.A1(_10198_),
    .A2(_03696_),
    .B1(_12044_),
    .B2(_10199_),
    .C1(_03166_),
    .C2(_10196_),
    .ZN(_10231_));
 AOI21_X2 _29183_ (.A(_10230_),
    .B1(_10231_),
    .B2(_10227_),
    .ZN(net204));
 CLKBUF_X3 _29184_ (.A(_03620_),
    .Z(_10232_));
 NOR2_X1 _29185_ (.A1(_10232_),
    .A2(net288),
    .ZN(_10233_));
 AOI222_X2 _29186_ (.A1(_10198_),
    .A2(_11158_),
    .B1(_12144_),
    .B2(_10199_),
    .C1(_03275_),
    .C2(_10196_),
    .ZN(_10234_));
 AOI21_X2 _29187_ (.A(_10233_),
    .B1(_10234_),
    .B2(_10227_),
    .ZN(net205));
 NOR2_X1 _29188_ (.A1(_10232_),
    .A2(net286),
    .ZN(_10235_));
 AOI222_X2 _29189_ (.A1(_10198_),
    .A2(_11202_),
    .B1(net327),
    .B2(_10199_),
    .C1(_03772_),
    .C2(_10196_),
    .ZN(_10236_));
 AOI21_X2 _29190_ (.A(_10235_),
    .B1(_10236_),
    .B2(_10227_),
    .ZN(net206));
 NAND2_X1 _29191_ (.A1(_10215_),
    .A2(_12316_),
    .ZN(_10237_));
 OAI221_X1 _29192_ (.A(_10237_),
    .B1(_11241_),
    .B2(_10217_),
    .C1(_10182_),
    .C2(_03660_),
    .ZN(_10238_));
 MUX2_X2 _29193_ (.A(_12985_),
    .B(_10238_),
    .S(_04153_),
    .Z(net207));
 NOR2_X1 _29194_ (.A1(_10232_),
    .A2(net292),
    .ZN(_10239_));
 AOI222_X2 _29195_ (.A1(_10197_),
    .A2(_03675_),
    .B1(_03727_),
    .B2(_10207_),
    .C1(_12392_),
    .C2(_10208_),
    .ZN(_10240_));
 AOI21_X4 _29196_ (.A(_10239_),
    .B1(_10240_),
    .B2(_10227_),
    .ZN(net208));
 NOR2_X1 _29197_ (.A1(_10232_),
    .A2(net314),
    .ZN(_10241_));
 AOI222_X2 _29198_ (.A1(_10197_),
    .A2(_10973_),
    .B1(_03736_),
    .B2(_10207_),
    .C1(net346),
    .C2(_10208_),
    .ZN(_10242_));
 AOI21_X2 _29199_ (.A(_10241_),
    .B1(_10242_),
    .B2(_10227_),
    .ZN(net209));
 NOR2_X1 _29200_ (.A1(_10232_),
    .A2(_13224_),
    .ZN(_10243_));
 AOI222_X2 _29201_ (.A1(_10197_),
    .A2(_11019_),
    .B1(_11351_),
    .B2(_10207_),
    .C1(net280),
    .C2(_10208_),
    .ZN(_10244_));
 AOI21_X2 _29202_ (.A(_10243_),
    .B1(_10244_),
    .B2(_10227_),
    .ZN(net210));
 NOR2_X1 _29203_ (.A1(_10232_),
    .A2(net330),
    .ZN(_10245_));
 BUF_X4 _29204_ (.A(_10196_),
    .Z(_10246_));
 AOI222_X2 _29205_ (.A1(_10246_),
    .A2(_03519_),
    .B1(net303),
    .B2(_10207_),
    .C1(_12651_),
    .C2(_10208_),
    .ZN(_10247_));
 AOI21_X4 _29206_ (.A(_10245_),
    .B1(_10247_),
    .B2(_10227_),
    .ZN(net211));
 NOR2_X1 _29207_ (.A1(_10232_),
    .A2(_03166_),
    .ZN(_10248_));
 AOI222_X2 _29208_ (.A1(_10246_),
    .A2(_03696_),
    .B1(_12044_),
    .B2(_10207_),
    .C1(net289),
    .C2(_10208_),
    .ZN(_10249_));
 AOI21_X4 _29209_ (.A(_10248_),
    .B1(_10249_),
    .B2(_10227_),
    .ZN(net212));
 AOI22_X1 _29210_ (.A1(_10189_),
    .A2(_12482_),
    .B1(net313),
    .B2(_10215_),
    .ZN(_10250_));
 OAI21_X1 _29211_ (.A(_10250_),
    .B1(_11313_),
    .B2(_10182_),
    .ZN(_10251_));
 MUX2_X2 _29212_ (.A(_10973_),
    .B(_10251_),
    .S(_04153_),
    .Z(net213));
 NOR2_X1 _29213_ (.A1(_10232_),
    .A2(_03275_),
    .ZN(_10252_));
 AOI222_X2 _29214_ (.A1(_10246_),
    .A2(_11158_),
    .B1(_12144_),
    .B2(_10207_),
    .C1(net287),
    .C2(_10215_),
    .ZN(_10253_));
 AOI21_X4 _29215_ (.A(_10252_),
    .B1(_10253_),
    .B2(_10194_),
    .ZN(net214));
 NOR2_X1 _29216_ (.A1(_10232_),
    .A2(_03772_),
    .ZN(_10254_));
 AOI222_X2 _29217_ (.A1(_10246_),
    .A2(_11202_),
    .B1(_12221_),
    .B2(_10189_),
    .C1(net285),
    .C2(_10215_),
    .ZN(_10255_));
 AOI21_X4 _29218_ (.A(_10254_),
    .B1(_10255_),
    .B2(_10194_),
    .ZN(net215));
 NOR2_X1 _29219_ (.A1(_10232_),
    .A2(_11019_),
    .ZN(_10256_));
 AOI222_X2 _29220_ (.A1(_10246_),
    .A2(_11351_),
    .B1(net280),
    .B2(_10189_),
    .C1(net329),
    .C2(_10215_),
    .ZN(_10257_));
 AOI21_X4 _29221_ (.A(_10256_),
    .B1(_10257_),
    .B2(_10194_),
    .ZN(net216));
 NOR2_X1 _29222_ (.A1(_04153_),
    .A2(_03519_),
    .ZN(_10258_));
 AOI222_X2 _29223_ (.A1(_10246_),
    .A2(net303),
    .B1(net355),
    .B2(_10189_),
    .C1(net330),
    .C2(_10215_),
    .ZN(_10259_));
 AOI21_X4 _29224_ (.A(_10258_),
    .B1(_10259_),
    .B2(_10194_),
    .ZN(net217));
 NOR2_X1 _29225_ (.A1(_04153_),
    .A2(_03696_),
    .ZN(_10260_));
 AOI222_X2 _29226_ (.A1(_10246_),
    .A2(_12044_),
    .B1(net289),
    .B2(_10189_),
    .C1(_03166_),
    .C2(_10215_),
    .ZN(_10261_));
 AOI21_X4 _29227_ (.A(_10260_),
    .B1(_10261_),
    .B2(_10194_),
    .ZN(net218));
 NOR2_X1 _29228_ (.A1(_04153_),
    .A2(_11158_),
    .ZN(_10262_));
 AOI222_X2 _29229_ (.A1(_10246_),
    .A2(_12144_),
    .B1(net287),
    .B2(_10189_),
    .C1(_03275_),
    .C2(_10215_),
    .ZN(_10263_));
 AOI21_X4 _29230_ (.A(_10262_),
    .B1(_10263_),
    .B2(_10194_),
    .ZN(net219));
 NOR2_X1 _29231_ (.A1(_04153_),
    .A2(_11202_),
    .ZN(_10264_));
 AOI222_X2 _29232_ (.A1(_10246_),
    .A2(_12221_),
    .B1(net285),
    .B2(_10189_),
    .C1(_03772_),
    .C2(_10215_),
    .ZN(_10265_));
 AOI21_X4 _29233_ (.A(_10264_),
    .B1(_10265_),
    .B2(_10194_),
    .ZN(net220));
 AOI22_X1 _29234_ (.A1(_07446_),
    .A2(_12316_),
    .B1(_12985_),
    .B2(_10188_),
    .ZN(_10266_));
 OAI21_X1 _29235_ (.A(_10266_),
    .B1(_03660_),
    .B2(_10216_),
    .ZN(_10267_));
 NOR2_X1 _29236_ (.A1(_03619_),
    .A2(_10267_),
    .ZN(_10268_));
 AOI21_X4 _29237_ (.A(_10268_),
    .B1(_11241_),
    .B2(_03619_),
    .ZN(net221));
 NOR2_X1 _29238_ (.A1(_04153_),
    .A2(_03727_),
    .ZN(_10269_));
 AOI222_X2 _29239_ (.A1(_10246_),
    .A2(net344),
    .B1(net292),
    .B2(_10189_),
    .C1(_10208_),
    .C2(_03675_),
    .ZN(_10270_));
 AOI21_X4 _29240_ (.A(_10269_),
    .B1(_10270_),
    .B2(_10194_),
    .ZN(net222));
 AND3_X1 _29241_ (.A1(_11418_),
    .A2(_03886_),
    .A3(_06323_),
    .ZN(\id_stage_i.branch_set_d ));
 NAND2_X1 _29242_ (.A1(net103),
    .A2(net254),
    .ZN(_10271_));
 NOR2_X1 _29243_ (.A1(_03960_),
    .A2(_10271_),
    .ZN(_10272_));
 OAI21_X1 _29244_ (.A(_04155_),
    .B1(net134),
    .B2(_03939_),
    .ZN(_10273_));
 AOI21_X1 _29245_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .B1(_03939_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_10274_));
 AOI22_X1 _29246_ (.A1(_07143_),
    .A2(_10273_),
    .B1(_10274_),
    .B2(_07144_),
    .ZN(_10275_));
 OR2_X1 _29247_ (.A1(_10272_),
    .A2(_10275_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NAND2_X1 _29248_ (.A1(_04155_),
    .A2(_10272_),
    .ZN(_10276_));
 AOI21_X1 _29249_ (.A(_07144_),
    .B1(_10274_),
    .B2(_10276_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 OR2_X1 _29250_ (.A1(_07156_),
    .A2(_07142_),
    .ZN(_10277_));
 NAND2_X1 _29251_ (.A1(_07150_),
    .A2(_07156_),
    .ZN(_10278_));
 AND3_X1 _29252_ (.A1(_07229_),
    .A2(_10277_),
    .A3(_10278_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 NOR2_X1 _29253_ (.A1(_06265_),
    .A2(_07155_),
    .ZN(_10279_));
 OAI21_X1 _29254_ (.A(_06858_),
    .B1(_10279_),
    .B2(_07142_),
    .ZN(_10280_));
 NOR2_X1 _29255_ (.A1(_07164_),
    .A2(_10280_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 NOR3_X1 _29256_ (.A1(_06893_),
    .A2(_10279_),
    .A3(_07162_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 NAND2_X1 _29257_ (.A1(_00134_),
    .A2(net134),
    .ZN(_10281_));
 NAND2_X1 _29258_ (.A1(_04155_),
    .A2(_10281_),
    .ZN(_10282_));
 NAND2_X1 _29259_ (.A1(_10271_),
    .A2(_10282_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 NAND3_X1 _29260_ (.A1(_04155_),
    .A2(net103),
    .A3(net254),
    .ZN(_10283_));
 AOI21_X1 _29261_ (.A(_07144_),
    .B1(_10283_),
    .B2(_00134_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AOI21_X1 _29262_ (.A(net103),
    .B1(_04162_),
    .B2(_00133_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 NAND2_X1 _29263_ (.A1(_03461_),
    .A2(_03854_),
    .ZN(_10284_));
 NAND4_X1 _29264_ (.A1(_10304_),
    .A2(_10284_),
    .A3(_03881_),
    .A4(_06287_),
    .ZN(_10285_));
 AOI21_X1 _29265_ (.A(_06265_),
    .B1(_06283_),
    .B2(_03931_),
    .ZN(_10286_));
 OAI22_X1 _29266_ (.A1(_06893_),
    .A2(_09783_),
    .B1(_10285_),
    .B2(_10286_),
    .ZN(\if_stage_i.instr_valid_id_d ));
 FA_X1 _29267_ (.A(_14065_),
    .B(_14064_),
    .CI(_14066_),
    .CO(_14067_),
    .S(_14068_));
 FA_X1 _29268_ (.A(_14069_),
    .B(_14070_),
    .CI(_14071_),
    .CO(_14072_),
    .S(_14073_));
 FA_X1 _29269_ (.A(_14074_),
    .B(_14075_),
    .CI(_14076_),
    .CO(_14077_),
    .S(_14078_));
 FA_X1 _29270_ (.A(_14079_),
    .B(_14080_),
    .CI(_14081_),
    .CO(_14082_),
    .S(_14083_));
 FA_X1 _29271_ (.A(_14084_),
    .B(_14085_),
    .CI(_14086_),
    .CO(_14087_),
    .S(_14088_));
 FA_X1 _29272_ (.A(_14089_),
    .B(_14090_),
    .CI(_14091_),
    .CO(_14092_),
    .S(_14093_));
 FA_X1 _29273_ (.A(_14094_),
    .B(_14095_),
    .CI(_14096_),
    .CO(_14097_),
    .S(_14098_));
 FA_X1 _29274_ (.A(_14099_),
    .B(_14100_),
    .CI(_14101_),
    .CO(_14102_),
    .S(_14103_));
 FA_X1 _29275_ (.A(_14104_),
    .B(_14105_),
    .CI(_14106_),
    .CO(_14107_),
    .S(_14108_));
 FA_X1 _29276_ (.A(_14109_),
    .B(_14110_),
    .CI(_14111_),
    .CO(_14112_),
    .S(_14113_));
 FA_X1 _29277_ (.A(_14092_),
    .B(_14114_),
    .CI(_14113_),
    .CO(_14115_),
    .S(_14116_));
 FA_X1 _29278_ (.A(_14117_),
    .B(_14118_),
    .CI(_14119_),
    .CO(_14120_),
    .S(_14121_));
 FA_X1 _29279_ (.A(_14122_),
    .B(_14123_),
    .CI(_14124_),
    .CO(_14125_),
    .S(_14126_));
 FA_X1 _29280_ (.A(_14127_),
    .B(_14128_),
    .CI(_14129_),
    .CO(_14130_),
    .S(_14131_));
 FA_X1 _29281_ (.A(_14132_),
    .B(_14133_),
    .CI(_14134_),
    .CO(_14135_),
    .S(_14136_));
 FA_X1 _29282_ (.A(_14112_),
    .B(_14137_),
    .CI(_14136_),
    .CO(_14138_),
    .S(_14139_));
 FA_X1 _29283_ (.A(_14140_),
    .B(_14141_),
    .CI(_14142_),
    .CO(_14143_),
    .S(_14144_));
 FA_X1 _29284_ (.A(_14145_),
    .B(_14146_),
    .CI(_14147_),
    .CO(_14148_),
    .S(_14149_));
 FA_X1 _29285_ (.A(_14150_),
    .B(_14151_),
    .CI(_14152_),
    .CO(_14153_),
    .S(_14154_));
 FA_X1 _29286_ (.A(_14155_),
    .B(_14156_),
    .CI(_14154_),
    .CO(_14157_),
    .S(_14158_));
 FA_X1 _29287_ (.A(_14159_),
    .B(_14160_),
    .CI(_14161_),
    .CO(_14162_),
    .S(_14163_));
 FA_X1 _29288_ (.A(_14164_),
    .B(_14163_),
    .CI(_14135_),
    .CO(_14165_),
    .S(_14166_));
 FA_X1 _29289_ (.A(_14167_),
    .B(_14168_),
    .CI(_14169_),
    .CO(_14170_),
    .S(_14171_));
 FA_X1 _29290_ (.A(_14172_),
    .B(_14173_),
    .CI(_14174_),
    .CO(_14175_),
    .S(_14176_));
 FA_X1 _29291_ (.A(_14177_),
    .B(_14178_),
    .CI(_14179_),
    .CO(_14180_),
    .S(_14181_));
 FA_X1 _29292_ (.A(_14182_),
    .B(_14183_),
    .CI(_14184_),
    .CO(_14185_),
    .S(_14186_));
 FA_X1 _29293_ (.A(_14187_),
    .B(_14181_),
    .CI(_14148_),
    .CO(_14188_),
    .S(_14189_));
 FA_X1 _29294_ (.A(_14190_),
    .B(_14191_),
    .CI(_14192_),
    .CO(_14193_),
    .S(_14194_));
 FA_X1 _29295_ (.A(_14195_),
    .B(_14194_),
    .CI(_14162_),
    .CO(_14196_),
    .S(_14197_));
 FA_X1 _29296_ (.A(_14198_),
    .B(_14199_),
    .CI(_14200_),
    .CO(_14201_),
    .S(_14202_));
 FA_X1 _29297_ (.A(_14203_),
    .B(_14204_),
    .CI(_14205_),
    .CO(_14206_),
    .S(_14207_));
 FA_X1 _29298_ (.A(_14208_),
    .B(_14210_),
    .CI(_14209_),
    .CO(_14211_),
    .S(_14212_));
 FA_X1 _29299_ (.A(_14213_),
    .B(_14214_),
    .CI(_14215_),
    .CO(_14216_),
    .S(_14217_));
 FA_X1 _29300_ (.A(_14212_),
    .B(_14180_),
    .CI(_14218_),
    .CO(_14219_),
    .S(_14220_));
 FA_X1 _29301_ (.A(_14221_),
    .B(_14222_),
    .CI(_14223_),
    .CO(_14224_),
    .S(_14225_));
 FA_X1 _29302_ (.A(_14226_),
    .B(_14225_),
    .CI(_14193_),
    .CO(_14227_),
    .S(_14228_));
 FA_X1 _29303_ (.A(_14229_),
    .B(_14230_),
    .CI(_14231_),
    .CO(_14232_),
    .S(_14233_));
 FA_X1 _29304_ (.A(_14234_),
    .B(_14235_),
    .CI(_14236_),
    .CO(_14237_),
    .S(_14238_));
 FA_X1 _29305_ (.A(_14239_),
    .B(_14240_),
    .CI(_14238_),
    .CO(_14241_),
    .S(_14242_));
 FA_X1 _29306_ (.A(_14243_),
    .B(_14244_),
    .CI(_14245_),
    .CO(_14246_),
    .S(_14247_));
 FA_X1 _29307_ (.A(_14248_),
    .B(_14250_),
    .CI(_14249_),
    .CO(_14251_),
    .S(_14252_));
 FA_X1 _29308_ (.A(_14253_),
    .B(_14254_),
    .CI(_14255_),
    .CO(_14256_),
    .S(_14257_));
 FA_X1 _29309_ (.A(_14252_),
    .B(_14211_),
    .CI(_14258_),
    .CO(_14259_),
    .S(_14260_));
 FA_X1 _29310_ (.A(_14261_),
    .B(_14262_),
    .CI(_14263_),
    .CO(_14264_),
    .S(_14265_));
 FA_X1 _29311_ (.A(_14266_),
    .B(_14224_),
    .CI(_14265_),
    .CO(_14267_),
    .S(_14268_));
 FA_X1 _29312_ (.A(_14269_),
    .B(_14270_),
    .CI(_14271_),
    .CO(_14272_),
    .S(_14273_));
 FA_X1 _29313_ (.A(_14274_),
    .B(_14275_),
    .CI(_14276_),
    .CO(_14277_),
    .S(_14278_));
 FA_X1 _29314_ (.A(_14279_),
    .B(_14232_),
    .CI(_14280_),
    .CO(_14281_),
    .S(_14282_));
 FA_X1 _29315_ (.A(_14283_),
    .B(_14284_),
    .CI(_14285_),
    .CO(_14286_),
    .S(_14287_));
 FA_X1 _29316_ (.A(_14288_),
    .B(_14290_),
    .CI(_14289_),
    .CO(_14291_),
    .S(_14292_));
 FA_X1 _29317_ (.A(_14293_),
    .B(_14294_),
    .CI(_14295_),
    .CO(_14296_),
    .S(_14297_));
 FA_X1 _29318_ (.A(_14298_),
    .B(_14251_),
    .CI(_14292_),
    .CO(_14299_),
    .S(_14300_));
 FA_X1 _29319_ (.A(_14301_),
    .B(_14259_),
    .CI(_14300_),
    .CO(_14302_),
    .S(_14303_));
 FA_X1 _29320_ (.A(_14305_),
    .B(_14304_),
    .CI(_14306_),
    .CO(_14307_),
    .S(_14308_));
 FA_X1 _29321_ (.A(_14309_),
    .B(_14308_),
    .CI(_14264_),
    .CO(_14310_),
    .S(_14311_));
 FA_X1 _29322_ (.A(_14312_),
    .B(_14313_),
    .CI(_14314_),
    .CO(_14315_),
    .S(_14316_));
 FA_X1 _29323_ (.A(_14317_),
    .B(_14319_),
    .CI(_14318_),
    .CO(_14320_),
    .S(_14321_));
 FA_X1 _29324_ (.A(_14322_),
    .B(_14272_),
    .CI(_14323_),
    .CO(_14324_),
    .S(_14325_));
 FA_X1 _29325_ (.A(_14326_),
    .B(_14327_),
    .CI(_14328_),
    .CO(_14329_),
    .S(_14330_));
 FA_X1 _29326_ (.A(_14331_),
    .B(_14333_),
    .CI(_14332_),
    .CO(_14334_),
    .S(_14335_));
 FA_X1 _29327_ (.A(_14336_),
    .B(_14337_),
    .CI(_14338_),
    .CO(_14339_),
    .S(_14340_));
 FA_X1 _29328_ (.A(_14341_),
    .B(_14291_),
    .CI(_14335_),
    .CO(_14342_),
    .S(_14343_));
 FA_X1 _29329_ (.A(_14344_),
    .B(_14299_),
    .CI(_14343_),
    .CO(_14345_),
    .S(_14346_));
 FA_X1 _29330_ (.A(_14347_),
    .B(_14348_),
    .CI(_14349_),
    .CO(_14350_),
    .S(_14351_));
 FA_X1 _29331_ (.A(_14352_),
    .B(_14353_),
    .CI(_14354_),
    .CO(_14355_),
    .S(_14356_));
 FA_X1 _29332_ (.A(_14357_),
    .B(_14356_),
    .CI(_14307_),
    .CO(_14358_),
    .S(_14359_));
 FA_X1 _29333_ (.A(_14360_),
    .B(_14361_),
    .CI(_14362_),
    .CO(_14363_),
    .S(_14364_));
 FA_X1 _29334_ (.A(_14351_),
    .B(_14364_),
    .CI(_14365_),
    .CO(_14366_),
    .S(_14367_));
 FA_X1 _29335_ (.A(_14368_),
    .B(_14369_),
    .CI(_14315_),
    .CO(_14370_),
    .S(_14371_));
 FA_X1 _29336_ (.A(_14372_),
    .B(_14373_),
    .CI(_14374_),
    .CO(_14375_),
    .S(_14376_));
 FA_X1 _29337_ (.A(_14377_),
    .B(_14378_),
    .CI(_14379_),
    .CO(_14380_),
    .S(_14381_));
 FA_X1 _29338_ (.A(_14381_),
    .B(_14329_),
    .CI(_14382_),
    .CO(_14383_),
    .S(_14384_));
 FA_X1 _29339_ (.A(_14385_),
    .B(_14386_),
    .CI(_14387_),
    .CO(_14388_),
    .S(_14389_));
 FA_X1 _29340_ (.A(_14390_),
    .B(_14391_),
    .CI(_14392_),
    .CO(_14393_),
    .S(_14394_));
 FA_X1 _29341_ (.A(_14395_),
    .B(_14334_),
    .CI(_14389_),
    .CO(_14396_),
    .S(_14397_));
 FA_X1 _29342_ (.A(_14398_),
    .B(_14342_),
    .CI(_14397_),
    .CO(_14399_),
    .S(_14400_));
 FA_X1 _29343_ (.A(_14401_),
    .B(_14402_),
    .CI(_14403_),
    .CO(_14404_),
    .S(_14405_));
 FA_X1 _29344_ (.A(_14406_),
    .B(_14407_),
    .CI(_14408_),
    .CO(_14409_),
    .S(_14410_));
 FA_X1 _29345_ (.A(_14411_),
    .B(_14410_),
    .CI(_14355_),
    .CO(_14412_),
    .S(_14413_));
 FA_X1 _29346_ (.A(_14414_),
    .B(_14415_),
    .CI(_14416_),
    .CO(_14417_),
    .S(_14418_));
 FA_X1 _29347_ (.A(_14421_),
    .B(_14420_),
    .CI(_14419_),
    .CO(_14422_),
    .S(_14423_));
 FA_X1 _29348_ (.A(_14423_),
    .B(_14424_),
    .CI(_14425_),
    .CO(_14426_),
    .S(_14427_));
 FA_X1 _29349_ (.A(_14428_),
    .B(_14429_),
    .CI(_14430_),
    .CO(_14431_),
    .S(_14432_));
 FA_X1 _29350_ (.A(_14433_),
    .B(_14434_),
    .CI(_14435_),
    .CO(_14436_),
    .S(_14437_));
 FA_X1 _29351_ (.A(_14437_),
    .B(_14380_),
    .CI(_14438_),
    .CO(_14439_),
    .S(_14440_));
 FA_X1 _29352_ (.A(_14441_),
    .B(_14442_),
    .CI(_14443_),
    .CO(_14444_),
    .S(_14445_));
 FA_X1 _29353_ (.A(_14446_),
    .B(_14447_),
    .CI(_14448_),
    .CO(_14449_),
    .S(_14450_));
 FA_X1 _29354_ (.A(_14451_),
    .B(_14388_),
    .CI(_14445_),
    .CO(_14452_),
    .S(_14453_));
 FA_X1 _29355_ (.A(_14383_),
    .B(_14453_),
    .CI(_14396_),
    .CO(_14454_),
    .S(_14455_));
 FA_X1 _29356_ (.A(_14457_),
    .B(_14456_),
    .CI(_14458_),
    .CO(_14459_),
    .S(_14460_));
 FA_X1 _29357_ (.A(_14461_),
    .B(_14462_),
    .CI(_14463_),
    .CO(_14464_),
    .S(_14465_));
 FA_X1 _29358_ (.A(_14466_),
    .B(_14465_),
    .CI(_14409_),
    .CO(_14467_),
    .S(_14468_));
 FA_X1 _29359_ (.A(_14469_),
    .B(_14470_),
    .CI(_14471_),
    .CO(_14472_),
    .S(_14473_));
 FA_X1 _29360_ (.A(_14476_),
    .B(_14474_),
    .CI(_14475_),
    .CO(_14477_),
    .S(_14478_));
 FA_X1 _29361_ (.A(_14479_),
    .B(_14478_),
    .CI(_14422_),
    .CO(_14480_),
    .S(_14481_));
 FA_X1 _29362_ (.A(_14482_),
    .B(_14483_),
    .CI(_14484_),
    .CO(_14485_),
    .S(_14486_));
 FA_X1 _29363_ (.A(_14489_),
    .B(_14488_),
    .CI(_14487_),
    .CO(_14490_),
    .S(_14491_));
 FA_X1 _29364_ (.A(_14431_),
    .B(_14491_),
    .CI(_14436_),
    .CO(_14492_),
    .S(_14493_));
 FA_X1 _29365_ (.A(_14494_),
    .B(_14495_),
    .CI(_14496_),
    .CO(_14497_),
    .S(_14498_));
 FA_X1 _29366_ (.A(_14499_),
    .B(_14501_),
    .CI(_14500_),
    .CO(_14502_),
    .S(_14503_));
 FA_X1 _29367_ (.A(_14504_),
    .B(_14505_),
    .CI(_14506_),
    .CO(_14507_),
    .S(_14508_));
 FA_X1 _29368_ (.A(_14509_),
    .B(_14444_),
    .CI(_14503_),
    .CO(_14510_),
    .S(_14511_));
 FA_X1 _29369_ (.A(_14439_),
    .B(_14452_),
    .CI(_14511_),
    .CO(_14512_),
    .S(_14513_));
 FA_X1 _29370_ (.A(_14514_),
    .B(_14515_),
    .CI(_14498_),
    .CO(_14516_),
    .S(_14517_));
 FA_X1 _29371_ (.A(_14518_),
    .B(_14519_),
    .CI(_14520_),
    .CO(_14521_),
    .S(_14522_));
 FA_X1 _29372_ (.A(_14523_),
    .B(_14522_),
    .CI(_14464_),
    .CO(_14524_),
    .S(_14525_));
 FA_X1 _29373_ (.A(_14526_),
    .B(_14527_),
    .CI(_14528_),
    .CO(_14529_),
    .S(_14530_));
 FA_X1 _29374_ (.A(_14533_),
    .B(_14532_),
    .CI(_14531_),
    .CO(_14534_),
    .S(_14535_));
 FA_X1 _29375_ (.A(_14536_),
    .B(_14477_),
    .CI(_14535_),
    .CO(_14537_),
    .S(_14538_));
 FA_X1 _29376_ (.A(_14539_),
    .B(_14540_),
    .CI(_14541_),
    .CO(_14542_),
    .S(_14543_));
 FA_X1 _29377_ (.A(_14544_),
    .B(_14545_),
    .CI(_14546_),
    .CO(_14547_),
    .S(_14548_));
 FA_X1 _29378_ (.A(_14550_),
    .B(_14548_),
    .CI(_14549_),
    .CO(_14551_),
    .S(_14552_));
 FA_X1 _29379_ (.A(_14553_),
    .B(_14555_),
    .CI(_14554_),
    .CO(_14556_),
    .S(_14557_));
 FA_X1 _29380_ (.A(_14557_),
    .B(_14490_),
    .CI(_14558_),
    .CO(_14559_),
    .S(_14560_));
 FA_X1 _29381_ (.A(_14552_),
    .B(_14561_),
    .CI(_14562_),
    .CO(_14563_),
    .S(_14564_));
 FA_X1 _29382_ (.A(_14565_),
    .B(_14566_),
    .CI(_14567_),
    .CO(_14568_),
    .S(_14569_));
 FA_X1 _29383_ (.A(_14570_),
    .B(_14571_),
    .CI(_14572_),
    .CO(_14573_),
    .S(_14574_));
 FA_X1 _29384_ (.A(_14569_),
    .B(_14502_),
    .CI(_14575_),
    .CO(_14576_),
    .S(_14577_));
 FA_X1 _29385_ (.A(_14492_),
    .B(_14577_),
    .CI(_14510_),
    .CO(_14578_),
    .S(_14579_));
 FA_X1 _29386_ (.A(_14580_),
    .B(_14581_),
    .CI(_14579_),
    .CO(_14582_),
    .S(_14583_));
 FA_X1 _29387_ (.A(_14584_),
    .B(_14585_),
    .CI(_14586_),
    .CO(_14587_),
    .S(_14588_));
 FA_X1 _29388_ (.A(_14589_),
    .B(_14521_),
    .CI(_14590_),
    .CO(_14591_),
    .S(_14592_));
 FA_X1 _29389_ (.A(net335),
    .B(_14594_),
    .CI(_14595_),
    .CO(_14596_),
    .S(_14597_));
 FA_X1 _29390_ (.A(_14598_),
    .B(_14597_),
    .CI(_14599_),
    .CO(_14600_),
    .S(_14601_));
 FA_X1 _29391_ (.A(_14603_),
    .B(_14602_),
    .CI(_14583_),
    .CO(_14604_),
    .S(_14605_));
 FA_X1 _29392_ (.A(_14605_),
    .B(_14534_),
    .CI(_14606_),
    .CO(_14607_),
    .S(_14608_));
 FA_X1 _29393_ (.A(_14609_),
    .B(_14610_),
    .CI(_14611_),
    .CO(_14612_),
    .S(_14613_));
 FA_X1 _29394_ (.A(_14614_),
    .B(_14615_),
    .CI(_14616_),
    .CO(_14617_),
    .S(_14618_));
 FA_X1 _29395_ (.A(_14619_),
    .B(_14613_),
    .CI(_14542_),
    .CO(_14620_),
    .S(_14621_));
 FA_X1 _29396_ (.A(_14622_),
    .B(_14623_),
    .CI(_14624_),
    .CO(_14625_),
    .S(_14626_));
 FA_X1 _29397_ (.A(_14627_),
    .B(_14626_),
    .CI(_14556_),
    .CO(_14628_),
    .S(_14629_));
 FA_X1 _29398_ (.A(_14630_),
    .B(_14629_),
    .CI(_14621_),
    .CO(_14631_),
    .S(_14632_));
 FA_X1 _29399_ (.A(_14633_),
    .B(_14634_),
    .CI(_14635_),
    .CO(_14636_),
    .S(_14637_));
 FA_X1 _29400_ (.A(_14638_),
    .B(_14639_),
    .CI(_14640_),
    .CO(_14641_),
    .S(_14642_));
 FA_X1 _29401_ (.A(_14643_),
    .B(_14637_),
    .CI(_14568_),
    .CO(_14644_),
    .S(_14645_));
 FA_X1 _29402_ (.A(_14559_),
    .B(_14645_),
    .CI(_14576_),
    .CO(_14646_),
    .S(_14647_));
 FA_X1 _29403_ (.A(_14632_),
    .B(_14648_),
    .CI(_14647_),
    .CO(_14649_),
    .S(_14650_));
 FA_X1 _29404_ (.A(_14651_),
    .B(_14586_),
    .CI(_14652_),
    .CO(_14653_),
    .S(_14654_));
 FA_X1 _29405_ (.A(_14655_),
    .B(_14656_),
    .CI(_14657_),
    .CO(_14658_),
    .S(_14659_));
 FA_X1 _29406_ (.A(_14660_),
    .B(_14661_),
    .CI(_14578_),
    .CO(_14662_),
    .S(_14663_));
 FA_X1 _29407_ (.A(_14650_),
    .B(_14582_),
    .CI(_14663_),
    .CO(_14664_),
    .S(_14665_));
 FA_X1 _29408_ (.A(_14665_),
    .B(_14604_),
    .CI(_14666_),
    .CO(_14667_),
    .S(_14668_));
 FA_X1 _29409_ (.A(_14669_),
    .B(_14670_),
    .CI(_14671_),
    .CO(_14672_),
    .S(_14673_));
 FA_X1 _29410_ (.A(_14674_),
    .B(_14675_),
    .CI(_14676_),
    .CO(_14677_),
    .S(_14678_));
 FA_X1 _29411_ (.A(_14612_),
    .B(_14679_),
    .CI(_14673_),
    .CO(_14680_),
    .S(_14681_));
 FA_X1 _29412_ (.A(_14682_),
    .B(_14683_),
    .CI(_14684_),
    .CO(_14685_),
    .S(_14686_));
 FA_X1 _29413_ (.A(_14686_),
    .B(_14625_),
    .CI(_14687_),
    .CO(_14688_),
    .S(_14689_));
 FA_X1 _29414_ (.A(_14689_),
    .B(_14681_),
    .CI(_14620_),
    .CO(_14690_),
    .S(_14691_));
 FA_X1 _29415_ (.A(_14692_),
    .B(_14693_),
    .CI(_14694_),
    .CO(_14695_),
    .S(_14696_));
 FA_X1 _29416_ (.A(_14697_),
    .B(_14698_),
    .CI(_14699_),
    .CO(_14700_),
    .S(_14701_));
 FA_X1 _29417_ (.A(_14636_),
    .B(_14702_),
    .CI(_14696_),
    .CO(_14703_),
    .S(_14704_));
 FA_X1 _29418_ (.A(_14628_),
    .B(_14704_),
    .CI(_14644_),
    .CO(_14705_),
    .S(_14706_));
 FA_X1 _29419_ (.A(_14631_),
    .B(_14706_),
    .CI(_14691_),
    .CO(_14707_),
    .S(_14708_));
 FA_X1 _29420_ (.A(_14651_),
    .B(_14709_),
    .CI(_14586_),
    .CO(_14710_),
    .S(_14711_));
 FA_X1 _29421_ (.A(_14712_),
    .B(_14713_),
    .CI(_14714_),
    .CO(_14715_),
    .S(_14716_));
 FA_X1 _29422_ (.A(_14717_),
    .B(_14718_),
    .CI(_14719_),
    .CO(_14720_),
    .S(_14721_));
 FA_X1 _29423_ (.A(_14649_),
    .B(_14722_),
    .CI(_14708_),
    .CO(_14723_),
    .S(_14724_));
 FA_X1 _29424_ (.A(_14724_),
    .B(_14664_),
    .CI(_14662_),
    .CO(_14725_),
    .S(_14726_));
 FA_X1 _29425_ (.A(_14727_),
    .B(_14728_),
    .CI(_14729_),
    .CO(_14730_),
    .S(_14731_));
 FA_X1 _29426_ (.A(_14732_),
    .B(_14733_),
    .CI(_14734_),
    .CO(_14735_),
    .S(_14736_));
 FA_X1 _29427_ (.A(_14672_),
    .B(_14737_),
    .CI(_14731_),
    .CO(_14738_),
    .S(_14739_));
 FA_X1 _29428_ (.A(_14740_),
    .B(_14741_),
    .CI(_14742_),
    .CO(_14743_),
    .S(_14744_));
 FA_X1 _29429_ (.A(_14744_),
    .B(_14685_),
    .CI(_14745_),
    .CO(_14746_),
    .S(_14747_));
 FA_X1 _29430_ (.A(_14747_),
    .B(_14739_),
    .CI(_14680_),
    .CO(_14748_),
    .S(_14749_));
 FA_X1 _29431_ (.A(_14750_),
    .B(_14751_),
    .CI(_14752_),
    .CO(_14753_),
    .S(_14754_));
 FA_X1 _29432_ (.A(_14755_),
    .B(_14756_),
    .CI(_14757_),
    .CO(_14758_),
    .S(_14759_));
 FA_X1 _29433_ (.A(_14695_),
    .B(_14754_),
    .CI(_14759_),
    .CO(_14760_),
    .S(_14761_));
 FA_X1 _29434_ (.A(_14688_),
    .B(_14761_),
    .CI(_14703_),
    .CO(_14762_),
    .S(_14763_));
 FA_X1 _29435_ (.A(_14690_),
    .B(_14763_),
    .CI(_14749_),
    .CO(_14764_),
    .S(_14765_));
 FA_X1 _29436_ (.A(_14651_),
    .B(_14586_),
    .CI(_14766_),
    .CO(_14767_),
    .S(_14768_));
 FA_X1 _29437_ (.A(_14769_),
    .B(_14770_),
    .CI(_14771_),
    .CO(_14772_),
    .S(_14773_));
 FA_X1 _29438_ (.A(_14774_),
    .B(_14775_),
    .CI(_14776_),
    .CO(_14777_),
    .S(_14778_));
 FA_X1 _29439_ (.A(_14765_),
    .B(_14707_),
    .CI(_14779_),
    .CO(_14780_),
    .S(_14781_));
 FA_X1 _29440_ (.A(_14781_),
    .B(_14723_),
    .CI(_14782_),
    .CO(_14783_),
    .S(_14784_));
 FA_X1 _29441_ (.A(_14785_),
    .B(_14786_),
    .CI(_14787_),
    .CO(_14788_),
    .S(_14789_));
 FA_X1 _29442_ (.A(_14790_),
    .B(_14791_),
    .CI(_14792_),
    .CO(_14793_),
    .S(_14794_));
 FA_X1 _29443_ (.A(_14795_),
    .B(_14789_),
    .CI(_14730_),
    .CO(_14796_),
    .S(_14797_));
 FA_X1 _29444_ (.A(_14798_),
    .B(_14799_),
    .CI(_14800_),
    .CO(_14801_),
    .S(_14802_));
 FA_X1 _29445_ (.A(_14803_),
    .B(_14802_),
    .CI(_14743_),
    .CO(_14804_),
    .S(_14805_));
 FA_X1 _29446_ (.A(_14738_),
    .B(_14805_),
    .CI(_14797_),
    .CO(_14806_),
    .S(_14807_));
 FA_X1 _29447_ (.A(_14808_),
    .B(_14809_),
    .CI(_14810_),
    .CO(_14811_),
    .S(_14812_));
 FA_X1 _29448_ (.A(_14813_),
    .B(_14814_),
    .CI(_14699_),
    .CO(_14815_),
    .S(_14816_));
 FA_X1 _29449_ (.A(_14812_),
    .B(_14753_),
    .CI(_14817_),
    .CO(_14818_),
    .S(_14819_));
 FA_X1 _29450_ (.A(_14819_),
    .B(_14760_),
    .CI(_14746_),
    .CO(_14820_),
    .S(_14821_));
 FA_X1 _29451_ (.A(_14821_),
    .B(_14807_),
    .CI(_14748_),
    .CO(_14822_),
    .S(_14823_));
 FA_X1 _29452_ (.A(_14651_),
    .B(_14824_),
    .CI(_14586_),
    .CO(_14825_),
    .S(_14826_));
 FA_X1 _29453_ (.A(_14827_),
    .B(_14758_),
    .CI(_14828_),
    .CO(_14829_),
    .S(_14830_));
 FA_X1 _29454_ (.A(_14831_),
    .B(_14832_),
    .CI(_14833_),
    .CO(_14834_),
    .S(_14835_));
 FA_X1 _29455_ (.A(_14764_),
    .B(_14836_),
    .CI(_14823_),
    .CO(_14837_),
    .S(_14838_));
 FA_X1 _29456_ (.A(_14780_),
    .B(_14839_),
    .CI(_14838_),
    .CO(_14840_),
    .S(_14841_));
 FA_X1 _29457_ (.A(_14842_),
    .B(_14843_),
    .CI(_14844_),
    .CO(_14845_),
    .S(_14846_));
 FA_X1 _29458_ (.A(_14847_),
    .B(_14848_),
    .CI(_14849_),
    .CO(_14850_),
    .S(_14851_));
 FA_X1 _29459_ (.A(_14846_),
    .B(_14788_),
    .CI(_14852_),
    .CO(_14853_),
    .S(_14854_));
 FA_X1 _29460_ (.A(_14855_),
    .B(_14856_),
    .CI(_14857_),
    .CO(_14858_),
    .S(_14859_));
 FA_X1 _29461_ (.A(_14859_),
    .B(_14801_),
    .CI(_14860_),
    .CO(_14861_),
    .S(_14862_));
 FA_X1 _29462_ (.A(_14862_),
    .B(_14854_),
    .CI(_14796_),
    .CO(_14863_),
    .S(_14864_));
 FA_X1 _29463_ (.A(_14865_),
    .B(_14866_),
    .CI(_14867_),
    .CO(_14868_),
    .S(_14869_));
 FA_X1 _29464_ (.A(_14869_),
    .B(_14811_),
    .CI(_14817_),
    .CO(_14870_),
    .S(_14871_));
 FA_X1 _29465_ (.A(_14804_),
    .B(_14871_),
    .CI(_14818_),
    .CO(_14872_),
    .S(_14873_));
 FA_X1 _29466_ (.A(_14864_),
    .B(_14806_),
    .CI(_14873_),
    .CO(_14874_),
    .S(_14875_));
 FA_X1 _29467_ (.A(_14651_),
    .B(net2),
    .CI(_14876_),
    .CO(_14877_),
    .S(_14878_));
 FA_X1 _29468_ (.A(_14879_),
    .B(_14880_),
    .CI(_14881_),
    .CO(_14882_),
    .S(_14883_));
 FA_X1 _29469_ (.A(_14884_),
    .B(_14885_),
    .CI(_14886_),
    .CO(_14887_),
    .S(_14888_));
 FA_X1 _29470_ (.A(_14875_),
    .B(_14822_),
    .CI(_14889_),
    .CO(_14890_),
    .S(_14891_));
 FA_X1 _29471_ (.A(_14891_),
    .B(_14837_),
    .CI(_14892_),
    .CO(_14893_),
    .S(_14894_));
 FA_X1 _29472_ (.A(_14895_),
    .B(_14896_),
    .CI(_14897_),
    .CO(_14898_),
    .S(_14899_));
 FA_X1 _29473_ (.A(_14900_),
    .B(_14901_),
    .CI(_14902_),
    .CO(_14903_),
    .S(_14904_));
 FA_X1 _29474_ (.A(_14845_),
    .B(_14905_),
    .CI(_14899_),
    .CO(_14906_),
    .S(_14907_));
 FA_X1 _29475_ (.A(_14908_),
    .B(_14909_),
    .CI(_14910_),
    .CO(_14911_),
    .S(_14912_));
 FA_X1 _29476_ (.A(_14912_),
    .B(_14858_),
    .CI(_14913_),
    .CO(_14914_),
    .S(_14915_));
 FA_X1 _29477_ (.A(_14915_),
    .B(_14907_),
    .CI(_14853_),
    .CO(_14916_),
    .S(_14917_));
 FA_X1 _29478_ (.A(_14866_),
    .B(_14918_),
    .CI(_14919_),
    .CO(_14920_),
    .S(_14921_));
 FA_X1 _29479_ (.A(_14922_),
    .B(_14816_),
    .CI(_14923_),
    .CO(_14924_),
    .S(_14925_));
 FA_X1 _29480_ (.A(_14861_),
    .B(_14926_),
    .CI(_14870_),
    .CO(_14927_),
    .S(_14928_));
 FA_X1 _29481_ (.A(_14863_),
    .B(_14928_),
    .CI(_14917_),
    .CO(_14929_),
    .S(_14930_));
 FA_X1 _29482_ (.A(_14651_),
    .B(_14931_),
    .CI(net2),
    .CO(_14932_),
    .S(_14933_));
 FA_X1 _29483_ (.A(_14934_),
    .B(_14935_),
    .CI(_14880_),
    .CO(_14936_),
    .S(_14937_));
 FA_X1 _29484_ (.A(_14938_),
    .B(_14939_),
    .CI(_14940_),
    .CO(_14941_),
    .S(_14942_));
 FA_X1 _29485_ (.A(_14930_),
    .B(_14943_),
    .CI(_14874_),
    .CO(_14944_),
    .S(_14945_));
 FA_X1 _29486_ (.A(_14890_),
    .B(_14946_),
    .CI(_14945_),
    .CO(_14947_),
    .S(_14948_));
 FA_X1 _29487_ (.A(_14949_),
    .B(_14950_),
    .CI(_14951_),
    .CO(_14952_),
    .S(_14953_));
 FA_X1 _29488_ (.A(_14954_),
    .B(_14955_),
    .CI(_14956_),
    .CO(_14957_),
    .S(_14958_));
 FA_X1 _29489_ (.A(_14958_),
    .B(_14953_),
    .CI(_14898_),
    .CO(_14959_),
    .S(_14960_));
 FA_X1 _29490_ (.A(_14961_),
    .B(_14962_),
    .CI(_14963_),
    .CO(_14964_),
    .S(_14965_));
 FA_X1 _29491_ (.A(_14966_),
    .B(_14965_),
    .CI(_14911_),
    .CO(_14967_),
    .S(_14968_));
 FA_X1 _29492_ (.A(_14906_),
    .B(_14968_),
    .CI(_14960_),
    .CO(_14969_),
    .S(_14970_));
 FA_X1 _29493_ (.A(_14971_),
    .B(_14972_),
    .CI(_14973_),
    .CO(_14974_),
    .S(_14975_));
 FA_X1 _29494_ (.A(_14817_),
    .B(_14976_),
    .CI(_14920_),
    .CO(_14977_),
    .S(_14978_));
 FA_X1 _29495_ (.A(_14978_),
    .B(_14979_),
    .CI(_14914_),
    .CO(_14980_),
    .S(_14981_));
 FA_X1 _29496_ (.A(_14981_),
    .B(_14970_),
    .CI(_14916_),
    .CO(_14982_),
    .S(_14983_));
 FA_X1 _29497_ (.A(_14984_),
    .B(_14651_),
    .CI(net2),
    .CO(_14985_),
    .S(_14986_));
 FA_X1 _29498_ (.A(_14987_),
    .B(_14880_),
    .CI(_14988_),
    .CO(_14989_),
    .S(_14990_));
 FA_X1 _29499_ (.A(_14991_),
    .B(_14992_),
    .CI(_14993_),
    .CO(_14994_),
    .S(_14995_));
 FA_X1 _29500_ (.A(_14929_),
    .B(_14983_),
    .CI(_14996_),
    .CO(_14997_),
    .S(_14998_));
 FA_X1 _29501_ (.A(_14998_),
    .B(_14944_),
    .CI(_14999_),
    .CO(_15000_),
    .S(_15001_));
 FA_X1 _29502_ (.A(_15002_),
    .B(_15003_),
    .CI(_15004_),
    .CO(_15005_),
    .S(_15006_));
 FA_X1 _29503_ (.A(_15007_),
    .B(_15008_),
    .CI(_15009_),
    .CO(_15010_),
    .S(_15011_));
 FA_X1 _29504_ (.A(_15006_),
    .B(_14952_),
    .CI(_15011_),
    .CO(_15012_),
    .S(_15013_));
 FA_X1 _29505_ (.A(_15014_),
    .B(_15015_),
    .CI(_15016_),
    .CO(_15017_),
    .S(_15018_));
 FA_X1 _29506_ (.A(_15018_),
    .B(_14964_),
    .CI(_14957_),
    .CO(_15019_),
    .S(_15020_));
 FA_X1 _29507_ (.A(_15020_),
    .B(_15013_),
    .CI(_14959_),
    .CO(_15021_),
    .S(_15022_));
 FA_X1 _29508_ (.A(_14816_),
    .B(_14975_),
    .CI(_14974_),
    .CO(_15023_),
    .S(_15024_));
 FA_X1 _29509_ (.A(_15025_),
    .B(_14977_),
    .CI(_14967_),
    .CO(_15026_),
    .S(_15027_));
 FA_X1 _29510_ (.A(_15022_),
    .B(_14969_),
    .CI(_15027_),
    .CO(_15028_),
    .S(_15029_));
 FA_X1 _29511_ (.A(_15030_),
    .B(_14651_),
    .CI(net1),
    .CO(_15031_),
    .S(_15032_));
 FA_X1 _29512_ (.A(_15033_),
    .B(_14880_),
    .CI(_15034_),
    .CO(_15035_),
    .S(_15036_));
 FA_X1 _29513_ (.A(_15037_),
    .B(_15038_),
    .CI(_15039_),
    .CO(_15040_),
    .S(_15041_));
 FA_X1 _29514_ (.A(_15042_),
    .B(_15029_),
    .CI(_14982_),
    .CO(_15043_),
    .S(_15044_));
 FA_X1 _29515_ (.A(_15044_),
    .B(_14997_),
    .CI(_15045_),
    .CO(_15046_),
    .S(_15047_));
 FA_X1 _29516_ (.A(_15048_),
    .B(_15049_),
    .CI(_15050_),
    .CO(_15051_),
    .S(_15052_));
 FA_X1 _29517_ (.A(_15053_),
    .B(_15054_),
    .CI(_15055_),
    .CO(_15056_),
    .S(_15057_));
 FA_X1 _29518_ (.A(_15052_),
    .B(_15057_),
    .CI(_15005_),
    .CO(_15058_),
    .S(_15059_));
 FA_X1 _29519_ (.A(_15060_),
    .B(_15061_),
    .CI(_15016_),
    .CO(_15062_),
    .S(_15063_));
 FA_X1 _29520_ (.A(_15017_),
    .B(_15010_),
    .CI(_15063_),
    .CO(_15064_),
    .S(_15065_));
 FA_X1 _29521_ (.A(_15059_),
    .B(_15012_),
    .CI(_15065_),
    .CO(_15066_),
    .S(_15067_));
 FA_X1 _29522_ (.A(_15025_),
    .B(_15019_),
    .CI(_15068_),
    .CO(_15069_),
    .S(_15070_));
 FA_X1 _29523_ (.A(_15021_),
    .B(_15070_),
    .CI(_15067_),
    .CO(_15071_),
    .S(_15072_));
 FA_X1 _29524_ (.A(_14651_),
    .B(net2),
    .CI(_15073_),
    .CO(_15074_),
    .S(_15075_));
 FA_X1 _29525_ (.A(_15076_),
    .B(_15077_),
    .CI(_14880_),
    .CO(_15078_),
    .S(_15079_));
 FA_X1 _29526_ (.A(_15080_),
    .B(_15081_),
    .CI(_15082_),
    .CO(_15083_),
    .S(_15084_));
 FA_X1 _29527_ (.A(_15072_),
    .B(_15085_),
    .CI(_15028_),
    .CO(_15086_),
    .S(_15087_));
 FA_X1 _29528_ (.A(_15087_),
    .B(_15043_),
    .CI(_15088_),
    .CO(_15089_),
    .S(_15090_));
 FA_X1 _29529_ (.A(_15091_),
    .B(_15092_),
    .CI(_15093_),
    .CO(_15094_),
    .S(_15095_));
 FA_X1 _29530_ (.A(_15096_),
    .B(_15097_),
    .CI(_15098_),
    .CO(_15099_),
    .S(_15100_));
 FA_X1 _29531_ (.A(_15100_),
    .B(_15051_),
    .CI(_15095_),
    .CO(_15101_),
    .S(_15102_));
 FA_X1 _29532_ (.A(_15103_),
    .B(_15104_),
    .CI(_15105_),
    .CO(_15106_),
    .S(_15107_));
 FA_X1 _29533_ (.A(_15062_),
    .B(_15056_),
    .CI(_15108_),
    .CO(_15109_),
    .S(_15110_));
 FA_X1 _29534_ (.A(_15058_),
    .B(_15102_),
    .CI(_15110_),
    .CO(_15111_),
    .S(_15112_));
 FA_X1 _29535_ (.A(_15025_),
    .B(_15064_),
    .CI(_15068_),
    .CO(_15113_),
    .S(_15114_));
 FA_X1 _29536_ (.A(_15066_),
    .B(_15112_),
    .CI(_15114_),
    .CO(_15115_),
    .S(_15116_));
 FA_X1 _29537_ (.A(_14651_),
    .B(_15117_),
    .CI(net1),
    .CO(_15118_),
    .S(_15119_));
 FA_X1 _29538_ (.A(_15120_),
    .B(_15121_),
    .CI(_14880_),
    .CO(_15122_),
    .S(_15123_));
 FA_X1 _29539_ (.A(_15124_),
    .B(_15125_),
    .CI(_15126_),
    .CO(_15127_),
    .S(_15128_));
 FA_X1 _29540_ (.A(_15071_),
    .B(_15116_),
    .CI(_15129_),
    .CO(_15130_),
    .S(_15131_));
 FA_X1 _29541_ (.A(_15086_),
    .B(_15132_),
    .CI(_15131_),
    .CO(_15133_),
    .S(_15134_));
 FA_X1 _29542_ (.A(_15135_),
    .B(_15136_),
    .CI(_15137_),
    .CO(_15138_),
    .S(_15139_));
 FA_X1 _29543_ (.A(_15140_),
    .B(_15141_),
    .CI(_15142_),
    .CO(_15143_),
    .S(_15144_));
 FA_X1 _29544_ (.A(_15139_),
    .B(_15144_),
    .CI(_15094_),
    .CO(_15145_),
    .S(_15146_));
 FA_X1 _29545_ (.A(_15099_),
    .B(_15147_),
    .CI(_15108_),
    .CO(_15148_),
    .S(_15149_));
 FA_X1 _29546_ (.A(_15149_),
    .B(_15146_),
    .CI(_15101_),
    .CO(_15150_),
    .S(_15151_));
 FA_X1 _29547_ (.A(_15025_),
    .B(_15068_),
    .CI(_15109_),
    .CO(_15152_),
    .S(_15153_));
 FA_X1 _29548_ (.A(_15153_),
    .B(_15111_),
    .CI(_15151_),
    .CO(_15154_),
    .S(_15155_));
 FA_X1 _29549_ (.A(_15156_),
    .B(_14651_),
    .CI(net1),
    .CO(_15157_),
    .S(_15158_));
 FA_X1 _29550_ (.A(_15159_),
    .B(_15160_),
    .CI(_14880_),
    .CO(_15161_),
    .S(_15162_));
 FA_X1 _29551_ (.A(_15163_),
    .B(_15164_),
    .CI(_15165_),
    .CO(_15166_),
    .S(_15167_));
 FA_X1 _29552_ (.A(_15168_),
    .B(_15115_),
    .CI(_15155_),
    .CO(_15169_),
    .S(_15170_));
 FA_X1 _29553_ (.A(_15130_),
    .B(_15171_),
    .CI(_15170_),
    .CO(_15172_),
    .S(_15173_));
 FA_X1 _29554_ (.A(_15174_),
    .B(_15175_),
    .CI(_15176_),
    .CO(_15177_),
    .S(_15178_));
 FA_X1 _29555_ (.A(_15179_),
    .B(_15180_),
    .CI(_15142_),
    .CO(_15181_),
    .S(_15182_));
 FA_X1 _29556_ (.A(_15178_),
    .B(_15182_),
    .CI(_15138_),
    .CO(_15183_),
    .S(_15184_));
 FA_X1 _29557_ (.A(_15147_),
    .B(_15143_),
    .CI(_15108_),
    .CO(_15185_),
    .S(_15186_));
 FA_X1 _29558_ (.A(_15184_),
    .B(_15145_),
    .CI(_15186_),
    .CO(_15187_),
    .S(_15188_));
 FA_X1 _29559_ (.A(_15025_),
    .B(_15068_),
    .CI(_15148_),
    .CO(_15189_),
    .S(_15190_));
 FA_X1 _29560_ (.A(_15190_),
    .B(_15188_),
    .CI(_15150_),
    .CO(_15191_),
    .S(_15192_));
 FA_X1 _29561_ (.A(_15193_),
    .B(_14651_),
    .CI(net1),
    .CO(_15194_),
    .S(_15195_));
 FA_X1 _29562_ (.A(_15196_),
    .B(_15197_),
    .CI(_14880_),
    .CO(_15198_),
    .S(_15199_));
 FA_X1 _29563_ (.A(_15200_),
    .B(_15201_),
    .CI(_15202_),
    .CO(_15203_),
    .S(_15204_));
 FA_X1 _29564_ (.A(_15192_),
    .B(_15205_),
    .CI(_15154_),
    .CO(_15206_),
    .S(_15207_));
 FA_X1 _29565_ (.A(_15169_),
    .B(_15208_),
    .CI(_15207_),
    .CO(_15209_),
    .S(_15210_));
 FA_X1 _29566_ (.A(_15211_),
    .B(_15212_),
    .CI(_15213_),
    .CO(_15214_),
    .S(_15215_));
 FA_X1 _29567_ (.A(_15216_),
    .B(_15217_),
    .CI(_15218_),
    .CO(_15219_),
    .S(_15220_));
 FA_X1 _29568_ (.A(_15215_),
    .B(_15177_),
    .CI(_15221_),
    .CO(_15222_),
    .S(_15223_));
 FA_X1 _29569_ (.A(_15147_),
    .B(_15181_),
    .CI(_15108_),
    .CO(_15224_),
    .S(_15225_));
 FA_X1 _29570_ (.A(_15223_),
    .B(_15183_),
    .CI(_15225_),
    .CO(_15226_),
    .S(_15227_));
 FA_X1 _29571_ (.A(_15025_),
    .B(_15185_),
    .CI(_15068_),
    .CO(_15228_),
    .S(_15229_));
 FA_X1 _29572_ (.A(_15227_),
    .B(_15187_),
    .CI(_15229_),
    .CO(_15230_),
    .S(_15231_));
 FA_X1 _29573_ (.A(_14651_),
    .B(net1),
    .CI(_15232_),
    .CO(_15233_),
    .S(_15234_));
 FA_X1 _29574_ (.A(_15235_),
    .B(_15236_),
    .CI(_14880_),
    .CO(_15237_),
    .S(_15238_));
 FA_X1 _29575_ (.A(_15239_),
    .B(_15240_),
    .CI(_15241_),
    .CO(_15242_),
    .S(_15243_));
 FA_X1 _29576_ (.A(_15231_),
    .B(_15244_),
    .CI(_15191_),
    .CO(_15245_),
    .S(_15246_));
 FA_X1 _29577_ (.A(_15246_),
    .B(_15206_),
    .CI(_15247_),
    .CO(_15248_),
    .S(_15249_));
 FA_X1 _29578_ (.A(_15250_),
    .B(_15251_),
    .CI(_15252_),
    .CO(_15253_),
    .S(_15254_));
 FA_X1 _29579_ (.A(_15220_),
    .B(_15255_),
    .CI(_15256_),
    .CO(_15257_),
    .S(_15258_));
 FA_X1 _29580_ (.A(_15147_),
    .B(_15259_),
    .CI(_15108_),
    .CO(_15260_),
    .S(_15261_));
 FA_X1 _29581_ (.A(_15262_),
    .B(_15222_),
    .CI(_15261_),
    .CO(_15263_),
    .S(_15264_));
 FA_X1 _29582_ (.A(_15024_),
    .B(_15266_),
    .CI(_15023_),
    .CO(_15267_),
    .S(_15268_));
 FA_X1 _29583_ (.A(_15264_),
    .B(_15226_),
    .CI(_15269_),
    .CO(_15270_),
    .S(_15271_));
 FA_X1 _29584_ (.A(_14651_),
    .B(_15272_),
    .CI(net1),
    .CO(_15273_),
    .S(_15274_));
 FA_X1 _29585_ (.A(_15275_),
    .B(_15276_),
    .CI(_14880_),
    .CO(_15277_),
    .S(_15278_));
 FA_X1 _29586_ (.A(_15279_),
    .B(_15280_),
    .CI(_15281_),
    .CO(_15282_),
    .S(_15283_));
 FA_X1 _29587_ (.A(_15271_),
    .B(_15230_),
    .CI(_15284_),
    .CO(_15285_),
    .S(_15286_));
 FA_X1 _29588_ (.A(_15286_),
    .B(_15245_),
    .CI(_15287_),
    .CO(_15288_),
    .S(_15289_));
 FA_X1 _29589_ (.A(_15251_),
    .B(_15290_),
    .CI(_15291_),
    .CO(_15292_),
    .S(_15293_));
 FA_X1 _29590_ (.A(_15294_),
    .B(_15295_),
    .CI(_15220_),
    .CO(_15296_),
    .S(_15297_));
 FA_X1 _29591_ (.A(_15261_),
    .B(_15298_),
    .CI(_15299_),
    .CO(_15300_),
    .S(_15301_));
 FA_X1 _29592_ (.A(_15024_),
    .B(_15302_),
    .CI(_15023_),
    .CO(_15303_),
    .S(_15304_));
 FA_X1 _29593_ (.A(_15301_),
    .B(_15263_),
    .CI(_15305_),
    .CO(_15306_),
    .S(_15307_));
 FA_X1 _29594_ (.A(_15308_),
    .B(_14651_),
    .CI(net1),
    .CO(_15309_),
    .S(_15310_));
 FA_X1 _29595_ (.A(_15311_),
    .B(_15312_),
    .CI(_14880_),
    .CO(_15313_),
    .S(_15314_));
 FA_X1 _29596_ (.A(_15315_),
    .B(_15316_),
    .CI(_15267_),
    .CO(_15317_),
    .S(_15318_));
 FA_X1 _29597_ (.A(_15307_),
    .B(_15270_),
    .CI(_15319_),
    .CO(_15320_),
    .S(_15321_));
 FA_X1 _29598_ (.A(_15322_),
    .B(_15321_),
    .CI(_15285_),
    .CO(_15323_),
    .S(_15324_));
 FA_X1 _29599_ (.A(_15251_),
    .B(_15325_),
    .CI(_15291_),
    .CO(_15326_),
    .S(_15327_));
 FA_X1 _29600_ (.A(_15220_),
    .B(_15328_),
    .CI(_15329_),
    .CO(_15330_),
    .S(_15331_));
 FA_X1 _29601_ (.A(_15331_),
    .B(_15296_),
    .CI(_15265_),
    .CO(_15332_),
    .S(_15333_));
 FA_X1 _29602_ (.A(_15334_),
    .B(_15300_),
    .CI(_15305_),
    .CO(_15335_),
    .S(_15336_));
 FA_X1 _29603_ (.A(_15337_),
    .B(_14651_),
    .CI(net1),
    .CO(_15338_),
    .S(_15339_));
 FA_X1 _29604_ (.A(_15339_),
    .B(_15309_),
    .CI(_14815_),
    .CO(_15340_),
    .S(_15341_));
 FA_X1 _29605_ (.A(_15342_),
    .B(_15303_),
    .CI(_15343_),
    .CO(_15344_),
    .S(_15345_));
 FA_X1 _29606_ (.A(_15346_),
    .B(_15336_),
    .CI(_15306_),
    .CO(_15347_),
    .S(_15348_));
 FA_X1 _29607_ (.A(_15349_),
    .B(_15348_),
    .CI(_15320_),
    .CO(_15350_),
    .S(_15351_));
 FA_X1 _29608_ (.A(_15352_),
    .B(_15353_),
    .CI(_15354_),
    .CO(_15355_),
    .S(_15356_));
 HA_X1 _29609_ (.A(_15357_),
    .B(_15358_),
    .CO(_15359_),
    .S(_15360_));
 HA_X1 _29610_ (.A(_15361_),
    .B(_15357_),
    .CO(_15362_),
    .S(_15363_));
 HA_X1 _29611_ (.A(_15364_),
    .B(_15358_),
    .CO(_15365_),
    .S(_15366_));
 HA_X1 _29612_ (.A(_15361_),
    .B(_15364_),
    .CO(_15367_),
    .S(_15368_));
 HA_X1 _29613_ (.A(_15369_),
    .B(_15370_),
    .CO(_15371_),
    .S(_15372_));
 HA_X1 _29614_ (.A(_14065_),
    .B(_14066_),
    .CO(_15373_),
    .S(_15374_));
 HA_X1 _29615_ (.A(_15375_),
    .B(_15376_),
    .CO(_15377_),
    .S(_15378_));
 HA_X1 _29616_ (.A(_15379_),
    .B(_15380_),
    .CO(_15381_),
    .S(_15382_));
 HA_X1 _29617_ (.A(_15383_),
    .B(_15384_),
    .CO(_15385_),
    .S(_15386_));
 HA_X1 _29618_ (.A(_15387_),
    .B(_15388_),
    .CO(_15389_),
    .S(_15390_));
 HA_X1 _29619_ (.A(_15391_),
    .B(_15392_),
    .CO(_15393_),
    .S(_15394_));
 HA_X1 _29620_ (.A(_15395_),
    .B(_15396_),
    .CO(_15397_),
    .S(_15398_));
 HA_X1 _29621_ (.A(_15399_),
    .B(_15400_),
    .CO(_15401_),
    .S(_15402_));
 HA_X1 _29622_ (.A(_15403_),
    .B(_15404_),
    .CO(_15405_),
    .S(_15406_));
 HA_X1 _29623_ (.A(_15407_),
    .B(_15408_),
    .CO(_15409_),
    .S(_15410_));
 HA_X1 _29624_ (.A(_15411_),
    .B(_15412_),
    .CO(_15413_),
    .S(_15414_));
 HA_X1 _29625_ (.A(_15415_),
    .B(_15416_),
    .CO(_15417_),
    .S(_15418_));
 HA_X1 _29626_ (.A(_15419_),
    .B(_15420_),
    .CO(_15421_),
    .S(_15422_));
 HA_X1 _29627_ (.A(_15423_),
    .B(_15424_),
    .CO(_15425_),
    .S(_15426_));
 HA_X1 _29628_ (.A(_15427_),
    .B(_15428_),
    .CO(_15429_),
    .S(_15430_));
 HA_X1 _29629_ (.A(_15431_),
    .B(_15432_),
    .CO(_15433_),
    .S(_15434_));
 HA_X1 _29630_ (.A(_15435_),
    .B(_15436_),
    .CO(_15437_),
    .S(_15438_));
 HA_X1 _29631_ (.A(_15439_),
    .B(_15440_),
    .CO(_15441_),
    .S(_15442_));
 HA_X1 _29632_ (.A(_15443_),
    .B(_15444_),
    .CO(_15445_),
    .S(_15446_));
 HA_X1 _29633_ (.A(_15447_),
    .B(_15448_),
    .CO(_15449_),
    .S(_15450_));
 HA_X1 _29634_ (.A(_15451_),
    .B(_15452_),
    .CO(_15453_),
    .S(_15454_));
 HA_X1 _29635_ (.A(_15455_),
    .B(_15456_),
    .CO(_15457_),
    .S(_15458_));
 HA_X1 _29636_ (.A(_15459_),
    .B(_15460_),
    .CO(_15461_),
    .S(_15462_));
 HA_X1 _29637_ (.A(_15463_),
    .B(_15464_),
    .CO(_15465_),
    .S(_15466_));
 HA_X1 _29638_ (.A(_15467_),
    .B(_15468_),
    .CO(_15469_),
    .S(_15470_));
 HA_X1 _29639_ (.A(_15471_),
    .B(_15472_),
    .CO(_15473_),
    .S(_15474_));
 HA_X1 _29640_ (.A(_15475_),
    .B(_15476_),
    .CO(_15477_),
    .S(_15478_));
 HA_X1 _29641_ (.A(_15479_),
    .B(_15480_),
    .CO(_15481_),
    .S(_15482_));
 HA_X1 _29642_ (.A(_15483_),
    .B(_15484_),
    .CO(_15485_),
    .S(_15486_));
 HA_X1 _29643_ (.A(_15487_),
    .B(_15488_),
    .CO(_15489_),
    .S(_15490_));
 HA_X1 _29644_ (.A(_15491_),
    .B(_15492_),
    .CO(_15493_),
    .S(_15494_));
 HA_X1 _29645_ (.A(_15495_),
    .B(_15496_),
    .CO(_15497_),
    .S(_15498_));
 HA_X1 _29646_ (.A(_15499_),
    .B(_15500_),
    .CO(_15501_),
    .S(_15502_));
 HA_X1 _29647_ (.A(_15503_),
    .B(\cs_registers_i.priv_lvl_q[0] ),
    .CO(_15504_),
    .S(_15505_));
 HA_X1 _29648_ (.A(_15506_),
    .B(_15507_),
    .CO(_15508_),
    .S(_15509_));
 HA_X1 _29649_ (.A(_15510_),
    .B(_15511_),
    .CO(_15512_),
    .S(_15513_));
 HA_X1 _29650_ (.A(_15510_),
    .B(_15514_),
    .CO(_15515_),
    .S(_15516_));
 HA_X1 _29651_ (.A(_15517_),
    .B(_15511_),
    .CO(_15518_),
    .S(_15519_));
 HA_X1 _29652_ (.A(_15517_),
    .B(_15514_),
    .CO(_15520_),
    .S(_15521_));
 HA_X1 _29653_ (.A(_15522_),
    .B(_15523_),
    .CO(_15524_),
    .S(_15525_));
 HA_X1 _29654_ (.A(_15522_),
    .B(_15526_),
    .CO(_15527_),
    .S(_15528_));
 HA_X1 _29655_ (.A(_15529_),
    .B(_15523_),
    .CO(_15530_),
    .S(_15531_));
 HA_X1 _29656_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .CO(_15532_),
    .S(_15533_));
 HA_X1 _29657_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .CO(_15534_),
    .S(_15535_));
 HA_X1 _29658_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CO(_15536_),
    .S(_15537_));
 HA_X1 _29659_ (.A(_15538_),
    .B(_15539_),
    .CO(_15540_),
    .S(_15541_));
 HA_X1 _29660_ (.A(_15538_),
    .B(_15539_),
    .CO(_15542_),
    .S(_15543_));
 HA_X1 _29661_ (.A(_15538_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_15544_),
    .S(_15545_));
 HA_X1 _29662_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_15539_),
    .CO(_15546_),
    .S(_15547_));
 HA_X1 _29663_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_15548_),
    .S(_15549_));
 HA_X1 _29664_ (.A(_15550_),
    .B(_15551_),
    .CO(_15552_),
    .S(_15553_));
 HA_X1 _29665_ (.A(_15552_),
    .B(_15554_),
    .CO(_15555_),
    .S(_15556_));
 HA_X1 _29666_ (.A(_15557_),
    .B(_15558_),
    .CO(_15559_),
    .S(_15560_));
 HA_X1 _29667_ (.A(_15555_),
    .B(_15560_),
    .CO(_15561_),
    .S(_15562_));
 HA_X1 _29668_ (.A(_15563_),
    .B(_15562_),
    .CO(_15564_),
    .S(_15565_));
 HA_X1 _29669_ (.A(_15566_),
    .B(_15567_),
    .CO(_14094_),
    .S(_15568_));
 HA_X1 _29670_ (.A(_15569_),
    .B(_15570_),
    .CO(_15571_),
    .S(_15572_));
 HA_X1 _29671_ (.A(_15572_),
    .B(_15559_),
    .CO(_15573_),
    .S(_15574_));
 HA_X1 _29672_ (.A(_15561_),
    .B(_15574_),
    .CO(_15575_),
    .S(_15576_));
 HA_X1 _29673_ (.A(_15568_),
    .B(_15576_),
    .CO(_15577_),
    .S(_15578_));
 HA_X1 _29674_ (.A(_15564_),
    .B(_15578_),
    .CO(_15579_),
    .S(_15580_));
 HA_X1 _29675_ (.A(_15571_),
    .B(_14098_),
    .CO(_15581_),
    .S(_15582_));
 HA_X1 _29676_ (.A(_15573_),
    .B(_15582_),
    .CO(_15583_),
    .S(_15584_));
 HA_X1 _29677_ (.A(_15584_),
    .B(_14088_),
    .CO(_15585_),
    .S(_15586_));
 HA_X1 _29678_ (.A(_15579_),
    .B(_15587_),
    .CO(_14124_),
    .S(_15588_));
 HA_X1 _29679_ (.A(_15589_),
    .B(_14108_),
    .CO(_15590_),
    .S(_15591_));
 HA_X1 _29680_ (.A(_15592_),
    .B(_14097_),
    .CO(_15593_),
    .S(_15594_));
 HA_X1 _29681_ (.A(_15581_),
    .B(_15594_),
    .CO(_15595_),
    .S(_15596_));
 HA_X1 _29682_ (.A(_15591_),
    .B(_15596_),
    .CO(_15597_),
    .S(_15598_));
 HA_X1 _29683_ (.A(_14122_),
    .B(_14123_),
    .CO(_15599_),
    .S(_15600_));
 HA_X1 _29684_ (.A(_15601_),
    .B(_15602_),
    .CO(_14155_),
    .S(_15603_));
 HA_X1 _29685_ (.A(_15603_),
    .B(_14131_),
    .CO(_15604_),
    .S(_15605_));
 HA_X1 _29686_ (.A(_15590_),
    .B(_15605_),
    .CO(_15606_),
    .S(_15607_));
 HA_X1 _29687_ (.A(_15608_),
    .B(_15609_),
    .CO(_15610_),
    .S(_15611_));
 HA_X1 _29688_ (.A(_15593_),
    .B(_15611_),
    .CO(_15612_),
    .S(_15613_));
 HA_X1 _29689_ (.A(_15613_),
    .B(_15607_),
    .CO(_15614_),
    .S(_15615_));
 HA_X1 _29690_ (.A(_15616_),
    .B(_15617_),
    .CO(_15618_),
    .S(_15619_));
 HA_X1 _29691_ (.A(_15604_),
    .B(_14158_),
    .CO(_15620_),
    .S(_15621_));
 HA_X1 _29692_ (.A(_15622_),
    .B(_15623_),
    .CO(_15624_),
    .S(_15625_));
 HA_X1 _29693_ (.A(_15621_),
    .B(_15626_),
    .CO(_14204_),
    .S(_15627_));
 HA_X1 _29694_ (.A(_15628_),
    .B(_15629_),
    .CO(_15630_),
    .S(_15631_));
 HA_X1 _29695_ (.A(_15632_),
    .B(_14157_),
    .CO(_15633_),
    .S(_15634_));
 HA_X1 _29696_ (.A(_15634_),
    .B(_15635_),
    .CO(_14236_),
    .S(_15636_));
 HA_X1 _29697_ (.A(_15637_),
    .B(_15638_),
    .CO(_15639_),
    .S(_15640_));
 HA_X1 _29698_ (.A(_15641_),
    .B(_15636_),
    .CO(_14239_),
    .S(_14203_));
 HA_X1 _29699_ (.A(_14207_),
    .B(_15642_),
    .CO(_15643_),
    .S(_15644_));
 HA_X1 _29700_ (.A(_15645_),
    .B(_15646_),
    .CO(_15647_),
    .S(_15648_));
 HA_X1 _29701_ (.A(_15649_),
    .B(_15650_),
    .CO(_15651_),
    .S(_15652_));
 HA_X1 _29702_ (.A(_15652_),
    .B(_15648_),
    .CO(_14276_),
    .S(_14234_));
 HA_X1 _29703_ (.A(_15653_),
    .B(_15654_),
    .CO(_15655_),
    .S(_15656_));
 HA_X1 _29704_ (.A(_14242_),
    .B(_14206_),
    .CO(_15657_),
    .S(_15658_));
 HA_X1 _29705_ (.A(_15659_),
    .B(_15647_),
    .CO(_15660_),
    .S(_15661_));
 HA_X1 _29706_ (.A(_15662_),
    .B(_15663_),
    .CO(_15664_),
    .S(_15665_));
 HA_X1 _29707_ (.A(_15665_),
    .B(_15661_),
    .CO(_14319_),
    .S(_14274_));
 HA_X1 _29708_ (.A(_15666_),
    .B(_15667_),
    .CO(_15668_),
    .S(_15669_));
 HA_X1 _29709_ (.A(_14241_),
    .B(_15670_),
    .CO(_15671_),
    .S(_15672_));
 HA_X1 _29710_ (.A(_15673_),
    .B(_15674_),
    .CO(_15675_),
    .S(_15676_));
 HA_X1 _29711_ (.A(_15676_),
    .B(_15677_),
    .CO(_14347_),
    .S(_15678_));
 HA_X1 _29712_ (.A(_15679_),
    .B(_15678_),
    .CO(_14365_),
    .S(_14317_));
 HA_X1 _29713_ (.A(_15681_),
    .B(_15680_),
    .CO(_14362_),
    .S(_15682_));
 HA_X1 _29714_ (.A(_15684_),
    .B(_15683_),
    .CO(_15685_),
    .S(_15686_));
 HA_X1 _29715_ (.A(_15687_),
    .B(_15688_),
    .CO(_15689_),
    .S(_15690_));
 HA_X1 _29716_ (.A(_15691_),
    .B(_15692_),
    .CO(_15693_),
    .S(_15694_));
 HA_X1 _29717_ (.A(_15690_),
    .B(_15694_),
    .CO(_14401_),
    .S(_14348_));
 HA_X1 _29718_ (.A(_15695_),
    .B(_15696_),
    .CO(_14416_),
    .S(_14360_));
 HA_X1 _29719_ (.A(_15698_),
    .B(_15697_),
    .CO(_15699_),
    .S(_15700_));
 HA_X1 _29720_ (.A(_14376_),
    .B(_15701_),
    .CO(_14456_),
    .S(_14402_));
 HA_X1 _29721_ (.A(_15702_),
    .B(_15703_),
    .CO(_14471_),
    .S(_14414_));
 HA_X1 _29722_ (.A(_15704_),
    .B(_15705_),
    .CO(_15706_),
    .S(_15707_));
 HA_X1 _29723_ (.A(_15708_),
    .B(_15709_),
    .CO(_14494_),
    .S(_15710_));
 HA_X1 _29724_ (.A(_15711_),
    .B(_15710_),
    .CO(_14514_),
    .S(_14458_));
 HA_X1 _29725_ (.A(_15712_),
    .B(_15713_),
    .CO(_14528_),
    .S(_14469_));
 HA_X1 _29726_ (.A(_15715_),
    .B(_15714_),
    .CO(_15716_),
    .S(_15717_));
 HA_X1 _29727_ (.A(_15718_),
    .B(_15719_),
    .CO(_14550_),
    .S(_15720_));
 HA_X1 _29728_ (.A(_15720_),
    .B(_14486_),
    .CO(_14562_),
    .S(_14495_));
 HA_X1 _29729_ (.A(_15721_),
    .B(_15722_),
    .CO(_14599_),
    .S(_14526_));
 HA_X1 _29730_ (.A(_15724_),
    .B(_15723_),
    .CO(_15725_),
    .S(_15726_));
 HA_X1 _29731_ (.A(_15728_),
    .B(_15727_),
    .CO(_15729_),
    .S(_15730_));
 HA_X1 _29732_ (.A(_14651_),
    .B(net1),
    .CO(_15731_),
    .S(_15732_));
 HA_X1 _29733_ (.A(_15733_),
    .B(_15734_),
    .CO(_14718_),
    .S(_15735_));
 HA_X1 _29734_ (.A(_15736_),
    .B(_15737_),
    .CO(_15738_),
    .S(_15739_));
 HA_X1 _29735_ (.A(_15740_),
    .B(_15741_),
    .CO(_14776_),
    .S(_14719_));
 HA_X1 _29736_ (.A(_15743_),
    .B(_15742_),
    .CO(_15744_),
    .S(_15745_));
 HA_X1 _29737_ (.A(_15746_),
    .B(_15747_),
    .CO(_14832_),
    .S(_14774_));
 HA_X1 _29738_ (.A(_15748_),
    .B(_15749_),
    .CO(_15750_),
    .S(_15751_));
 HA_X1 _29739_ (.A(_15752_),
    .B(_15753_),
    .CO(_14886_),
    .S(_14833_));
 HA_X1 _29740_ (.A(_15754_),
    .B(_15755_),
    .CO(_15756_),
    .S(_15757_));
 HA_X1 _29741_ (.A(_15758_),
    .B(_15759_),
    .CO(_14939_),
    .S(_14884_));
 HA_X1 _29742_ (.A(_15760_),
    .B(_15761_),
    .CO(_15762_),
    .S(_15763_));
 HA_X1 _29743_ (.A(_15764_),
    .B(_15765_),
    .CO(_14992_),
    .S(_14940_));
 HA_X1 _29744_ (.A(_15766_),
    .B(_15767_),
    .CO(_15768_),
    .S(_15769_));
 HA_X1 _29745_ (.A(_15770_),
    .B(_15771_),
    .CO(_15038_),
    .S(_14993_));
 HA_X1 _29746_ (.A(_15772_),
    .B(_15773_),
    .CO(_15774_),
    .S(_15775_));
 HA_X1 _29747_ (.A(_15776_),
    .B(_15777_),
    .CO(_15080_),
    .S(_15037_));
 HA_X1 _29748_ (.A(_15778_),
    .B(_15779_),
    .CO(_15780_),
    .S(_15781_));
 HA_X1 _29749_ (.A(_15782_),
    .B(_15783_),
    .CO(_15124_),
    .S(_15082_));
 HA_X1 _29750_ (.A(_15784_),
    .B(_15785_),
    .CO(_15786_),
    .S(_15787_));
 HA_X1 _29751_ (.A(_15788_),
    .B(_15789_),
    .CO(_15164_),
    .S(_15126_));
 HA_X1 _29752_ (.A(_15790_),
    .B(_15791_),
    .CO(_15792_),
    .S(_15793_));
 HA_X1 _29753_ (.A(_15794_),
    .B(_15795_),
    .CO(_15201_),
    .S(_15165_));
 HA_X1 _29754_ (.A(_15796_),
    .B(_15797_),
    .CO(_15798_),
    .S(_15799_));
 HA_X1 _29755_ (.A(_15800_),
    .B(_15801_),
    .CO(_15241_),
    .S(_15202_));
 HA_X1 _29756_ (.A(_15802_),
    .B(_15803_),
    .CO(_15804_),
    .S(_15805_));
 HA_X1 _29757_ (.A(_15806_),
    .B(_15807_),
    .CO(_15281_),
    .S(_15239_));
 HA_X1 _29758_ (.A(_15808_),
    .B(_15809_),
    .CO(_15810_),
    .S(_15811_));
 HA_X1 _29759_ (.A(_15812_),
    .B(_15813_),
    .CO(_15316_),
    .S(_15280_));
 HA_X1 _29760_ (.A(_15814_),
    .B(_15815_),
    .CO(_15816_),
    .S(_15817_));
 HA_X1 _29761_ (.A(_15818_),
    .B(_15819_),
    .CO(_15343_),
    .S(_15315_));
 HA_X1 _29762_ (.A(_15820_),
    .B(_15821_),
    .CO(_15822_),
    .S(_15823_));
 HA_X1 _29763_ (.A(_15824_),
    .B(_15825_),
    .CO(_15826_),
    .S(_15342_));
 HA_X1 _29764_ (.A(_15827_),
    .B(_15828_),
    .CO(_15829_),
    .S(_15830_));
 HA_X1 _29765_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_15831_),
    .CO(_15832_),
    .S(_15833_));
 HA_X1 _29766_ (.A(_15834_),
    .B(_15835_),
    .CO(_15836_),
    .S(_15837_));
 HA_X1 _29767_ (.A(_15835_),
    .B(_15838_),
    .CO(_15839_),
    .S(_15840_));
 HA_X1 _29768_ (.A(_15841_),
    .B(_15842_),
    .CO(_15843_),
    .S(_15844_));
 HA_X1 _29769_ (.A(_15845_),
    .B(_15846_),
    .CO(_15847_),
    .S(_15848_));
 HA_X1 _29770_ (.A(_15849_),
    .B(_15834_),
    .CO(_15850_),
    .S(_15851_));
 HA_X1 _29771_ (.A(_15852_),
    .B(_15853_),
    .CO(_15854_),
    .S(_15855_));
 HA_X1 _29772_ (.A(_15856_),
    .B(_15857_),
    .CO(_15858_),
    .S(_15859_));
 HA_X1 _29773_ (.A(_15860_),
    .B(_15861_),
    .CO(_15862_),
    .S(_15863_));
 HA_X1 _29774_ (.A(_15864_),
    .B(_15865_),
    .CO(_15866_),
    .S(_15867_));
 HA_X1 _29775_ (.A(_15868_),
    .B(_15869_),
    .CO(_15870_),
    .S(_15871_));
 HA_X1 _29776_ (.A(_15872_),
    .B(_15873_),
    .CO(_15874_),
    .S(_15875_));
 HA_X1 _29777_ (.A(_15876_),
    .B(_15877_),
    .CO(_15878_),
    .S(_15879_));
 HA_X1 _29778_ (.A(_15880_),
    .B(_15881_),
    .CO(_15882_),
    .S(_15883_));
 HA_X1 _29779_ (.A(_15884_),
    .B(_15885_),
    .CO(_15886_),
    .S(_15887_));
 HA_X1 _29780_ (.A(_15888_),
    .B(_15889_),
    .CO(_15890_),
    .S(_15891_));
 HA_X1 _29781_ (.A(_15892_),
    .B(_15893_),
    .CO(_15894_),
    .S(_15895_));
 HA_X1 _29782_ (.A(_15896_),
    .B(_15897_),
    .CO(_15898_),
    .S(_15899_));
 HA_X1 _29783_ (.A(_15900_),
    .B(_15901_),
    .CO(_15902_),
    .S(_15903_));
 HA_X1 _29784_ (.A(_15904_),
    .B(_15905_),
    .CO(_15906_),
    .S(_15907_));
 HA_X1 _29785_ (.A(_15908_),
    .B(_15909_),
    .CO(_15910_),
    .S(_15911_));
 HA_X1 _29786_ (.A(_15912_),
    .B(_15913_),
    .CO(_15914_),
    .S(_15915_));
 HA_X1 _29787_ (.A(_15916_),
    .B(_15917_),
    .CO(_15918_),
    .S(_15919_));
 HA_X1 _29788_ (.A(_15920_),
    .B(_15921_),
    .CO(_15922_),
    .S(_15923_));
 HA_X1 _29789_ (.A(_15924_),
    .B(_15925_),
    .CO(_15926_),
    .S(_15927_));
 HA_X1 _29790_ (.A(_15928_),
    .B(_15929_),
    .CO(_15930_),
    .S(_15931_));
 HA_X1 _29791_ (.A(_15932_),
    .B(_15933_),
    .CO(_15934_),
    .S(_15935_));
 HA_X1 _29792_ (.A(_15936_),
    .B(_15937_),
    .CO(_15938_),
    .S(_15939_));
 HA_X1 _29793_ (.A(_15940_),
    .B(_15941_),
    .CO(_15942_),
    .S(_15943_));
 HA_X1 _29794_ (.A(_15944_),
    .B(_15945_),
    .CO(_15946_),
    .S(_15947_));
 HA_X1 _29795_ (.A(_15948_),
    .B(_15949_),
    .CO(_15950_),
    .S(_15951_));
 HA_X1 _29796_ (.A(_15952_),
    .B(_15953_),
    .CO(_15954_),
    .S(_15955_));
 HA_X1 _29797_ (.A(_15956_),
    .B(_15957_),
    .CO(_15958_),
    .S(_15959_));
 HA_X1 _29798_ (.A(_15960_),
    .B(_15961_),
    .CO(_15962_),
    .S(_15963_));
 HA_X1 _29799_ (.A(_15964_),
    .B(_15965_),
    .CO(_15966_),
    .S(_15967_));
 HA_X1 _29800_ (.A(_15968_),
    .B(_15969_),
    .CO(_15970_),
    .S(_15971_));
 HA_X1 _29801_ (.A(_15972_),
    .B(_15973_),
    .CO(_15974_),
    .S(_15975_));
 HA_X1 _29802_ (.A(_15976_),
    .B(_15977_),
    .CO(_15978_),
    .S(_15979_));
 HA_X1 _29803_ (.A(_15980_),
    .B(_15981_),
    .CO(_15982_),
    .S(_15983_));
 HA_X1 _29804_ (.A(_15984_),
    .B(_15985_),
    .CO(_15986_),
    .S(_15987_));
 HA_X1 _29805_ (.A(_15988_),
    .B(_15989_),
    .CO(_15990_),
    .S(_15991_));
 HA_X1 _29806_ (.A(_15992_),
    .B(_15993_),
    .CO(_15994_),
    .S(_15995_));
 HA_X1 _29807_ (.A(_15996_),
    .B(_15997_),
    .CO(_15998_),
    .S(_15999_));
 HA_X1 _29808_ (.A(_16000_),
    .B(_16001_),
    .CO(_16002_),
    .S(_16003_));
 HA_X1 _29809_ (.A(_16004_),
    .B(_16005_),
    .CO(_16006_),
    .S(_16007_));
 HA_X1 _29810_ (.A(_16008_),
    .B(_16009_),
    .CO(_16010_),
    .S(_16011_));
 HA_X1 _29811_ (.A(_16012_),
    .B(_16013_),
    .CO(_16014_),
    .S(_16015_));
 HA_X1 _29812_ (.A(_16016_),
    .B(_16017_),
    .CO(_16018_),
    .S(_16019_));
 HA_X1 _29813_ (.A(_16020_),
    .B(_16021_),
    .CO(_16022_),
    .S(_16023_));
 HA_X1 _29814_ (.A(_16024_),
    .B(_16025_),
    .CO(_16026_),
    .S(_16027_));
 HA_X1 _29815_ (.A(_16028_),
    .B(_16029_),
    .CO(_16030_),
    .S(_16031_));
 HA_X1 _29816_ (.A(_16032_),
    .B(_16033_),
    .CO(_16034_),
    .S(_16035_));
 HA_X1 _29817_ (.A(_16036_),
    .B(_16037_),
    .CO(_16038_),
    .S(_16039_));
 HA_X1 _29818_ (.A(_16040_),
    .B(_16041_),
    .CO(_16042_),
    .S(_16043_));
 HA_X1 _29819_ (.A(_16044_),
    .B(_16045_),
    .CO(_16046_),
    .S(_16047_));
 HA_X1 _29820_ (.A(_16048_),
    .B(_16049_),
    .CO(_16050_),
    .S(_16051_));
 HA_X1 _29821_ (.A(_16052_),
    .B(_16053_),
    .CO(_16054_),
    .S(_16055_));
 HA_X1 _29822_ (.A(_16056_),
    .B(_16057_),
    .CO(_16058_),
    .S(_16059_));
 HA_X1 _29823_ (.A(_16060_),
    .B(_16061_),
    .CO(_16062_),
    .S(_16063_));
 HA_X1 _29824_ (.A(_16064_),
    .B(_16065_),
    .CO(_16066_),
    .S(_16067_));
 HA_X1 _29825_ (.A(_16068_),
    .B(_16069_),
    .CO(_16070_),
    .S(_16071_));
 HA_X1 _29826_ (.A(_16072_),
    .B(_16073_),
    .CO(_16074_),
    .S(_16075_));
 HA_X1 _29827_ (.A(_16076_),
    .B(_16077_),
    .CO(_16078_),
    .S(_16079_));
 HA_X1 _29828_ (.A(_16080_),
    .B(_16081_),
    .CO(_16082_),
    .S(_16083_));
 HA_X1 _29829_ (.A(_16084_),
    .B(_16085_),
    .CO(_16086_),
    .S(_16087_));
 HA_X1 _29830_ (.A(net15),
    .B(_16085_),
    .CO(_16088_),
    .S(_16089_));
 HA_X1 _29831_ (.A(_16090_),
    .B(_16085_),
    .CO(_16091_),
    .S(_16092_));
 HA_X1 _29832_ (.A(net15),
    .B(\alu_adder_result_ex[0] ),
    .CO(_16093_),
    .S(_16094_));
 HA_X1 _29833_ (.A(net15),
    .B(\alu_adder_result_ex[0] ),
    .CO(_16095_),
    .S(_16096_));
 HA_X1 _29834_ (.A(net15),
    .B(_14068_),
    .CO(_16097_),
    .S(_16098_));
 HA_X1 _29835_ (.A(net15),
    .B(_14068_),
    .CO(_16099_),
    .S(_16100_));
 HA_X1 _29836_ (.A(_16090_),
    .B(\alu_adder_result_ex[0] ),
    .CO(_16101_),
    .S(_16102_));
 HA_X1 _29837_ (.A(_16090_),
    .B(\alu_adder_result_ex[0] ),
    .CO(_16103_),
    .S(_16104_));
 HA_X1 _29838_ (.A(_16090_),
    .B(_14068_),
    .CO(_16105_),
    .S(_16106_));
 HA_X1 _29839_ (.A(_16107_),
    .B(_16108_),
    .CO(_16109_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 HA_X1 _29840_ (.A(_16109_),
    .B(_16110_),
    .CO(_16111_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 DFFR_X1 _29841_ (.D(_01680_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.data_type_q[2] ),
    .QN(_14049_));
 DFFR_X1 _29842_ (.D(_01681_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.data_type_q[1] ),
    .QN(_14048_));
 DFFR_X2 _29843_ (.D(_01682_),
    .RN(net263),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .QN(_14047_));
 DFFR_X1 _29844_ (.D(_01683_),
    .RN(net264),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .QN(_14046_));
 DFFR_X2 _29845_ (.D(_01684_),
    .RN(net264),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .QN(_00179_));
 DFFR_X1 _29846_ (.D(_01685_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .QN(_14045_));
 DFFS_X1 _29847_ (.D(_01686_),
    .SN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .QN(_14050_));
 CLKBUF_X3 clkbuf_regs_0_core_clock (.A(clk_i),
    .Z(delaynet_0_core_clock));
 BUF_X1 _29849_ (.A(net266),
    .Z(alert_major_o));
 BUF_X1 _29850_ (.A(net267),
    .Z(alert_minor_o));
 BUF_X1 _29851_ (.A(net268),
    .Z(data_addr_o[0]));
 BUF_X1 _29852_ (.A(net269),
    .Z(data_addr_o[1]));
 BUF_X2 _29853_ (.A(\alu_adder_result_ex[2] ),
    .Z(net176));
 BUF_X2 _29854_ (.A(\alu_adder_result_ex[3] ),
    .Z(net179));
 CLKBUF_X2 _29855_ (.A(\alu_adder_result_ex[4] ),
    .Z(net180));
 BUF_X2 _29856_ (.A(\alu_adder_result_ex[5] ),
    .Z(net181));
 BUF_X2 _29857_ (.A(\alu_adder_result_ex[6] ),
    .Z(net182));
 BUF_X1 _29858_ (.A(\alu_adder_result_ex[7] ),
    .Z(net183));
 CLKBUF_X2 _29859_ (.A(\alu_adder_result_ex[8] ),
    .Z(net184));
 BUF_X1 _29860_ (.A(\alu_adder_result_ex[9] ),
    .Z(net185));
 BUF_X1 _29861_ (.A(\alu_adder_result_ex[10] ),
    .Z(net156));
 BUF_X1 _29862_ (.A(\alu_adder_result_ex[11] ),
    .Z(net157));
 BUF_X2 _29863_ (.A(\alu_adder_result_ex[12] ),
    .Z(net158));
 BUF_X1 _29864_ (.A(\alu_adder_result_ex[13] ),
    .Z(net159));
 CLKBUF_X2 _29865_ (.A(\alu_adder_result_ex[14] ),
    .Z(net160));
 BUF_X1 _29866_ (.A(\alu_adder_result_ex[15] ),
    .Z(net161));
 BUF_X1 _29867_ (.A(\alu_adder_result_ex[16] ),
    .Z(net162));
 BUF_X1 _29868_ (.A(\alu_adder_result_ex[17] ),
    .Z(net163));
 BUF_X1 _29869_ (.A(net369),
    .Z(net164));
 BUF_X1 _29870_ (.A(\alu_adder_result_ex[19] ),
    .Z(net165));
 CLKBUF_X2 _29871_ (.A(\alu_adder_result_ex[20] ),
    .Z(net166));
 CLKBUF_X2 _29872_ (.A(\alu_adder_result_ex[21] ),
    .Z(net167));
 BUF_X2 _29873_ (.A(\alu_adder_result_ex[22] ),
    .Z(net168));
 BUF_X1 _29874_ (.A(net413),
    .Z(net169));
 CLKBUF_X2 _29875_ (.A(\alu_adder_result_ex[24] ),
    .Z(net170));
 BUF_X1 _29876_ (.A(\alu_adder_result_ex[25] ),
    .Z(net171));
 BUF_X1 _29877_ (.A(net382),
    .Z(net172));
 CLKBUF_X2 _29878_ (.A(net375),
    .Z(net173));
 CLKBUF_X2 _29879_ (.A(\alu_adder_result_ex[28] ),
    .Z(net174));
 BUF_X1 _29880_ (.A(\alu_adder_result_ex[29] ),
    .Z(net175));
 BUF_X2 _29881_ (.A(\alu_adder_result_ex[30] ),
    .Z(net177));
 BUF_X2 _29882_ (.A(\alu_adder_result_ex[31] ),
    .Z(net178));
 BUF_X1 _29883_ (.A(net270),
    .Z(instr_addr_o[0]));
 BUF_X1 _29884_ (.A(net271),
    .Z(instr_addr_o[1]));
 DFFR_X1 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .RN(net261),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(core_busy_q),
    .QN(_14044_));
 DLL_X1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00006_),
    .GN(clknet_leaf_107_clk_i_regs),
    .Q(\core_clock_gate_i.en_latch ));
 DFFR_X1 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_01687_),
    .RN(net262),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mcountinhibit[0] ),
    .QN(_00553_));
 DFFR_X2 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_01688_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mcountinhibit[2] ),
    .QN(_01159_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_01689_),
    .RN(net261),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .QN(_00551_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_01690_),
    .RN(net261),
    .CK(clknet_leaf_118_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .QN(_14043_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_01691_),
    .RN(net261),
    .CK(clknet_leaf_118_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .QN(_14042_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_01692_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .QN(_14041_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_01693_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .QN(_14040_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_01694_),
    .RN(net261),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .QN(_14039_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_01695_),
    .RN(net261),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .QN(_14038_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_01696_),
    .RN(net261),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .QN(_14037_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_01697_),
    .RN(net261),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .QN(_14036_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_01698_),
    .RN(net261),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .QN(_14035_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_01699_),
    .RN(net153),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .QN(_14034_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_01700_),
    .RN(net261),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .QN(_14033_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_01701_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .QN(_14032_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_01702_),
    .RN(net261),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .QN(_14031_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_01703_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .QN(_14030_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_01704_),
    .RN(net153),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .QN(_14029_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_01705_),
    .RN(net261),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .QN(_14028_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_01706_),
    .RN(net261),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .QN(_14027_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_01707_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .QN(_14026_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_01708_),
    .RN(net261),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .QN(_14025_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_01709_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .QN(_14024_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_01710_),
    .RN(net261),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .QN(_14023_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_01711_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .QN(_14022_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_01712_),
    .RN(net261),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .QN(_14021_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_01713_),
    .RN(net153),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .QN(_14020_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_01714_),
    .RN(net153),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .QN(_14019_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_01715_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .QN(_14018_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_01716_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .QN(_14017_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_01717_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .QN(_14016_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_01718_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .QN(_14015_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_01719_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .QN(_14014_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_01720_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .QN(_14013_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_01721_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .QN(_14012_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_01722_),
    .RN(net261),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .QN(_14011_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_01723_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .QN(_14010_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_01724_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .QN(_14009_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_01725_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .QN(_14008_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_01726_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .QN(_14007_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_01727_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .QN(_14006_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_01728_),
    .RN(net153),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .QN(_14005_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_01729_),
    .RN(net153),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .QN(_14004_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_01730_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .QN(_14003_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_01731_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .QN(_14002_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_01732_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .QN(_14001_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_01733_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .QN(_14000_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_01734_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .QN(_13999_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_01735_),
    .RN(net153),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .QN(_13998_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_01736_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .QN(_13997_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_01737_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .QN(_13996_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_01738_),
    .RN(net153),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .QN(_13995_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_01739_),
    .RN(net153),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .QN(_13994_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_01740_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .QN(_13993_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_01741_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .QN(_13992_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_01742_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .QN(_13991_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_01743_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .QN(_13990_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_01744_),
    .RN(net261),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .QN(_13989_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_01745_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .QN(_13988_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_01746_),
    .RN(net153),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .QN(_13987_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_01747_),
    .RN(net153),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .QN(_13986_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_01748_),
    .RN(net153),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .QN(_13985_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_01749_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .QN(_13984_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_01750_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .QN(_13983_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_01751_),
    .RN(net261),
    .CK(clknet_leaf_118_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .QN(_13982_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_01752_),
    .RN(net261),
    .CK(clknet_leaf_118_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .QN(_13981_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_01753_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mhpmcounter[2][0] ),
    .QN(_00552_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_01754_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][10] ),
    .QN(_13980_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_01755_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][11] ),
    .QN(_13979_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_01756_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][12] ),
    .QN(_13978_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_01757_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][13] ),
    .QN(_13977_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_01758_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][14] ),
    .QN(_13976_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_01759_),
    .RN(net261),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][15] ),
    .QN(_13975_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_01760_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][16] ),
    .QN(_13974_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_01761_),
    .RN(net261),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mhpmcounter[2][17] ),
    .QN(_13973_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_01762_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][18] ),
    .QN(_13972_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_01763_),
    .RN(net261),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[2][19] ),
    .QN(_13971_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_01764_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mhpmcounter[2][1] ),
    .QN(_13970_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_01765_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][20] ),
    .QN(_13969_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_01766_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][21] ),
    .QN(_13968_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_01767_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][22] ),
    .QN(_13967_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_01768_),
    .RN(net261),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mhpmcounter[2][23] ),
    .QN(_13966_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_01769_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][24] ),
    .QN(_13965_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_01770_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][25] ),
    .QN(_13964_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_01771_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][26] ),
    .QN(_13963_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_01772_),
    .RN(net261),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[2][27] ),
    .QN(_13962_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_01773_),
    .RN(net261),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mhpmcounter[2][28] ),
    .QN(_13961_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_01774_),
    .RN(net262),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mhpmcounter[2][29] ),
    .QN(_13960_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_01775_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][2] ),
    .QN(_13959_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_01776_),
    .RN(net261),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][30] ),
    .QN(_13958_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_01777_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][31] ),
    .QN(_13957_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_01778_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][32] ),
    .QN(_13956_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_01779_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][33] ),
    .QN(_13955_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_01780_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mhpmcounter[2][34] ),
    .QN(_13954_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_01781_),
    .RN(net261),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][35] ),
    .QN(_13953_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_01782_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.mhpmcounter[2][36] ),
    .QN(_13952_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_01783_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.mhpmcounter[2][37] ),
    .QN(_13951_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_01784_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][38] ),
    .QN(_13950_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_01785_),
    .RN(net261),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.mhpmcounter[2][39] ),
    .QN(_13949_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_01786_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mhpmcounter[2][3] ),
    .QN(_13948_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_01787_),
    .RN(net153),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][40] ),
    .QN(_13947_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_01788_),
    .RN(net153),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][41] ),
    .QN(_13946_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_01789_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mhpmcounter[2][42] ),
    .QN(_13945_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_01790_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mhpmcounter[2][43] ),
    .QN(_13944_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_01791_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mhpmcounter[2][44] ),
    .QN(_13943_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_01792_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mhpmcounter[2][45] ),
    .QN(_13942_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_01793_),
    .RN(net153),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][46] ),
    .QN(_13941_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_01794_),
    .RN(net153),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][47] ),
    .QN(_13940_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_01795_),
    .RN(net153),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.mhpmcounter[2][48] ),
    .QN(_13939_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_01796_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][49] ),
    .QN(_13938_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_01797_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][4] ),
    .QN(_13937_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_01798_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][50] ),
    .QN(_13936_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_01799_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][51] ),
    .QN(_13935_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_01800_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][52] ),
    .QN(_13934_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_01801_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][53] ),
    .QN(_13933_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_01802_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][54] ),
    .QN(_13932_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_01803_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][55] ),
    .QN(_13931_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_01804_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][56] ),
    .QN(_13930_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_01805_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][57] ),
    .QN(_13929_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_01806_),
    .RN(net153),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mhpmcounter[2][58] ),
    .QN(_13928_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_01807_),
    .RN(net153),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[2][59] ),
    .QN(_13927_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_01808_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][5] ),
    .QN(_13926_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_01809_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][60] ),
    .QN(_13925_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_01810_),
    .RN(net153),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[2][61] ),
    .QN(_13924_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_01811_),
    .RN(net153),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[2][62] ),
    .QN(_13923_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_01812_),
    .RN(net153),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[2][63] ),
    .QN(_13922_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_01813_),
    .RN(net261),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mhpmcounter[2][6] ),
    .QN(_13921_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_01814_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][7] ),
    .QN(_13920_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_01815_),
    .RN(net261),
    .CK(clknet_leaf_118_clk),
    .Q(\cs_registers_i.mhpmcounter[2][8] ),
    .QN(_13919_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_01816_),
    .RN(net261),
    .CK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mhpmcounter[2][9] ),
    .QN(_13918_));
 DFFS_X1 \cs_registers_i.priv_lvl_q[0]$_DFFE_PN1P_  (.D(_01817_),
    .SN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.priv_lvl_q[0] ),
    .QN(_13917_));
 DFFS_X1 \cs_registers_i.priv_lvl_q[1]$_DFFE_PN1P_  (.D(_01818_),
    .SN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.priv_lvl_q[1] ),
    .QN(_15500_));
 DFFS_X2 \cs_registers_i.u_dcsr_csr.rdata_q[0]$_DFFE_PN1P_  (.D(_01819_),
    .SN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[0] ),
    .QN(_13916_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01820_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.dcsr_q[11] ),
    .QN(_13915_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01821_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.dcsr_q[12] ),
    .QN(_13914_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01822_),
    .RN(net265),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.dcsr_q[13] ),
    .QN(_13913_));
 DFFR_X2 \cs_registers_i.u_dcsr_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01823_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.dcsr_q[15] ),
    .QN(_13912_));
 DFFS_X2 \cs_registers_i.u_dcsr_csr.rdata_q[1]$_DFFE_PN1P_  (.D(_01824_),
    .SN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.dcsr_q[1] ),
    .QN(_13911_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01825_),
    .RN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[2] ),
    .QN(_01162_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01826_),
    .RN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[6] ),
    .QN(_13910_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01827_),
    .RN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[7] ),
    .QN(_13909_));
 DFFR_X2 \cs_registers_i.u_dcsr_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01828_),
    .RN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.dcsr_q[8] ),
    .QN(_13908_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01829_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_depc_o[10] ),
    .QN(_13907_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01830_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.csr_depc_o[11] ),
    .QN(_13906_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01831_),
    .RN(net265),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_depc_o[12] ),
    .QN(_13905_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01832_),
    .RN(net265),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_depc_o[13] ),
    .QN(_13904_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01833_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_depc_o[14] ),
    .QN(_13903_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01834_),
    .RN(net264),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_depc_o[15] ),
    .QN(_13902_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01835_),
    .RN(net265),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.csr_depc_o[16] ),
    .QN(_13901_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01836_),
    .RN(net265),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_depc_o[17] ),
    .QN(_13900_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01837_),
    .RN(net265),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_depc_o[18] ),
    .QN(_13899_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01838_),
    .RN(net264),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_depc_o[19] ),
    .QN(_13898_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01839_),
    .RN(net262),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.csr_depc_o[1] ),
    .QN(_00554_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01840_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_depc_o[20] ),
    .QN(_13897_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01841_),
    .RN(net265),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_depc_o[21] ),
    .QN(_13896_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01842_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_depc_o[22] ),
    .QN(_13895_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01843_),
    .RN(net265),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_depc_o[23] ),
    .QN(_13894_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01844_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_depc_o[24] ),
    .QN(_13893_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01845_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_depc_o[25] ),
    .QN(_13892_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01846_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_depc_o[26] ),
    .QN(_13891_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01847_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_depc_o[27] ),
    .QN(_13890_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_01848_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_depc_o[28] ),
    .QN(_13889_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_01849_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_depc_o[29] ),
    .QN(_13888_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01850_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.csr_depc_o[2] ),
    .QN(_13887_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_01851_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_depc_o[30] ),
    .QN(_13886_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_01852_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_depc_o[31] ),
    .QN(_13885_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01853_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.csr_depc_o[3] ),
    .QN(_01163_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01854_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.csr_depc_o[4] ),
    .QN(_01164_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01855_),
    .RN(net265),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_depc_o[5] ),
    .QN(_01165_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01856_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.csr_depc_o[6] ),
    .QN(_01166_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01857_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.csr_depc_o[7] ),
    .QN(_13884_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01858_),
    .RN(net264),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_depc_o[8] ),
    .QN(_13883_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01859_),
    .RN(net265),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_depc_o[9] ),
    .QN(_13882_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01860_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.dscratch0_q[0] ),
    .QN(_13881_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01861_),
    .RN(net262),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.dscratch0_q[10] ),
    .QN(_13880_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01862_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.dscratch0_q[11] ),
    .QN(_13879_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01863_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.dscratch0_q[12] ),
    .QN(_13878_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01864_),
    .RN(net265),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.dscratch0_q[13] ),
    .QN(_13877_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01865_),
    .RN(net265),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.dscratch0_q[14] ),
    .QN(_13876_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01866_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.dscratch0_q[15] ),
    .QN(_13875_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01867_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.dscratch0_q[16] ),
    .QN(_13874_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01868_),
    .RN(net262),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch0_q[17] ),
    .QN(_13873_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01869_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.dscratch0_q[18] ),
    .QN(_13872_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01870_),
    .RN(net262),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.dscratch0_q[19] ),
    .QN(_13871_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01871_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch0_q[1] ),
    .QN(_13870_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01872_),
    .RN(net153),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.dscratch0_q[20] ),
    .QN(_13869_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01873_),
    .RN(net265),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.dscratch0_q[21] ),
    .QN(_13868_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01874_),
    .RN(net153),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.dscratch0_q[22] ),
    .QN(_13867_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01875_),
    .RN(net265),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.dscratch0_q[23] ),
    .QN(_13866_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01876_),
    .RN(net265),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.dscratch0_q[24] ),
    .QN(_13865_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01877_),
    .RN(net265),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.dscratch0_q[25] ),
    .QN(_13864_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01878_),
    .RN(net265),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.dscratch0_q[26] ),
    .QN(_13863_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01879_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch0_q[27] ),
    .QN(_13862_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_01880_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.dscratch0_q[28] ),
    .QN(_13861_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_01881_),
    .RN(net153),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.dscratch0_q[29] ),
    .QN(_13860_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01882_),
    .RN(net262),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.dscratch0_q[2] ),
    .QN(_13859_));
 DFFR_X2 \cs_registers_i.u_dscratch0_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_01883_),
    .RN(net153),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.dscratch0_q[30] ),
    .QN(_13858_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_01884_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch0_q[31] ),
    .QN(_13857_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01885_),
    .RN(net261),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch0_q[3] ),
    .QN(_13856_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01886_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch0_q[4] ),
    .QN(_13855_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01887_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[5] ),
    .QN(_13854_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01888_),
    .RN(net261),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch0_q[6] ),
    .QN(_13853_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01889_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[7] ),
    .QN(_13852_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01890_),
    .RN(net262),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch0_q[8] ),
    .QN(_13851_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01891_),
    .RN(net262),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.dscratch0_q[9] ),
    .QN(_13850_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01892_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.dscratch1_q[0] ),
    .QN(_13849_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01893_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[10] ),
    .QN(_13848_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01894_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.dscratch1_q[11] ),
    .QN(_13847_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01895_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.dscratch1_q[12] ),
    .QN(_13846_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01896_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch1_q[13] ),
    .QN(_13845_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01897_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.dscratch1_q[14] ),
    .QN(_13844_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01898_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch1_q[15] ),
    .QN(_13843_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01899_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.dscratch1_q[16] ),
    .QN(_13842_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01900_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.dscratch1_q[17] ),
    .QN(_13841_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01901_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.dscratch1_q[18] ),
    .QN(_13840_));
 DFFR_X2 \cs_registers_i.u_dscratch1_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01902_),
    .RN(net153),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.dscratch1_q[19] ),
    .QN(_13839_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01903_),
    .RN(net153),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch1_q[1] ),
    .QN(_13838_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01904_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[20] ),
    .QN(_13837_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01905_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch1_q[21] ),
    .QN(_13836_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01906_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[22] ),
    .QN(_13835_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01907_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.dscratch1_q[23] ),
    .QN(_13834_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01908_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.dscratch1_q[24] ),
    .QN(_13833_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01909_),
    .RN(net153),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.dscratch1_q[25] ),
    .QN(_13832_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01910_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[26] ),
    .QN(_13831_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01911_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[27] ),
    .QN(_13830_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_01912_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.dscratch1_q[28] ),
    .QN(_13829_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_01913_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[29] ),
    .QN(_13828_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01914_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch1_q[2] ),
    .QN(_13827_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_01915_),
    .RN(net153),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.dscratch1_q[30] ),
    .QN(_13826_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_01916_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.dscratch1_q[31] ),
    .QN(_13825_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01917_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[3] ),
    .QN(_13824_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01918_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch1_q[4] ),
    .QN(_13823_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01919_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[5] ),
    .QN(_13822_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01920_),
    .RN(net261),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.dscratch1_q[6] ),
    .QN(_13821_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01921_),
    .RN(net262),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[7] ),
    .QN(_13820_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01922_),
    .RN(net262),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch1_q[8] ),
    .QN(_13819_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01923_),
    .RN(net153),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.dscratch1_q[9] ),
    .QN(_13818_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01924_),
    .RN(net262),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mcause_q[0] ),
    .QN(_13817_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01925_),
    .RN(net262),
    .CK(clknet_leaf_57_clk),
    .Q(\cs_registers_i.mcause_q[1] ),
    .QN(_13816_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01926_),
    .RN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mcause_q[2] ),
    .QN(_13815_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01927_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mcause_q[3] ),
    .QN(_13814_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01928_),
    .RN(net265),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mcause_q[4] ),
    .QN(_13813_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01929_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mcause_q[5] ),
    .QN(_13812_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01930_),
    .RN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_mepc_o[0] ),
    .QN(_13811_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01931_),
    .RN(net265),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_mepc_o[10] ),
    .QN(_13810_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01932_),
    .RN(net264),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.csr_mepc_o[11] ),
    .QN(_13809_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01933_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_mepc_o[12] ),
    .QN(_13808_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01934_),
    .RN(net265),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.csr_mepc_o[13] ),
    .QN(_13807_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01935_),
    .RN(net153),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.csr_mepc_o[14] ),
    .QN(_13806_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01936_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.csr_mepc_o[15] ),
    .QN(_13805_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01937_),
    .RN(net153),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.csr_mepc_o[16] ),
    .QN(_13804_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01938_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.csr_mepc_o[17] ),
    .QN(_13803_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01939_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_mepc_o[18] ),
    .QN(_13802_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01940_),
    .RN(net265),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.csr_mepc_o[19] ),
    .QN(_13801_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01941_),
    .RN(net265),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.csr_mepc_o[1] ),
    .QN(_13800_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01942_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.csr_mepc_o[20] ),
    .QN(_13799_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01943_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.csr_mepc_o[21] ),
    .QN(_13798_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01944_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mepc_o[22] ),
    .QN(_13797_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01945_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.csr_mepc_o[23] ),
    .QN(_13796_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01946_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.csr_mepc_o[24] ),
    .QN(_13795_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01947_),
    .RN(net153),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.csr_mepc_o[25] ),
    .QN(_13794_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01948_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mepc_o[26] ),
    .QN(_13793_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01949_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_mepc_o[27] ),
    .QN(_13792_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_01950_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_mepc_o[28] ),
    .QN(_13791_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_01951_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_mepc_o[29] ),
    .QN(_13790_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01952_),
    .RN(net265),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.csr_mepc_o[2] ),
    .QN(_13789_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_01953_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_mepc_o[30] ),
    .QN(_13788_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_01954_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mepc_o[31] ),
    .QN(_13787_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01955_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.csr_mepc_o[3] ),
    .QN(_13786_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01956_),
    .RN(net265),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.csr_mepc_o[4] ),
    .QN(_13785_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01957_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mepc_o[5] ),
    .QN(_13784_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01958_),
    .RN(net264),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.csr_mepc_o[6] ),
    .QN(_13783_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01959_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.csr_mepc_o[7] ),
    .QN(_13782_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01960_),
    .RN(net264),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.csr_mepc_o[8] ),
    .QN(_13781_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01961_),
    .RN(net264),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.csr_mepc_o[9] ),
    .QN(_13780_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01962_),
    .RN(net265),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mie_q[0] ),
    .QN(_13779_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01963_),
    .RN(net153),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mie_q[10] ),
    .QN(_13778_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01964_),
    .RN(net265),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mie_q[11] ),
    .QN(_13777_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01965_),
    .RN(net153),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mie_q[12] ),
    .QN(_13776_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01966_),
    .RN(net153),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mie_q[13] ),
    .QN(_13775_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01967_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mie_q[14] ),
    .QN(_13774_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01968_),
    .RN(net262),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.mie_q[15] ),
    .QN(_13773_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01969_),
    .RN(net261),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.mie_q[16] ),
    .QN(_13772_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01970_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.mie_q[17] ),
    .QN(_13771_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01971_),
    .RN(net265),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mie_q[1] ),
    .QN(_13770_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_01972_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.mie_q[2] ),
    .QN(_13769_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_01973_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mie_q[3] ),
    .QN(_13768_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_01974_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mie_q[4] ),
    .QN(_13767_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_01975_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mie_q[5] ),
    .QN(_13766_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_01976_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mie_q[6] ),
    .QN(_13765_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_01977_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mie_q[7] ),
    .QN(_13764_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01978_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mie_q[8] ),
    .QN(_13763_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01979_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mie_q[9] ),
    .QN(_13762_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_01980_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[0] ),
    .QN(_13761_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_01981_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[10] ),
    .QN(_13760_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01982_),
    .RN(net265),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mscratch_q[11] ),
    .QN(_13759_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01983_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.mscratch_q[12] ),
    .QN(_13758_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01984_),
    .RN(net265),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.mscratch_q[13] ),
    .QN(_13757_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01985_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.mscratch_q[14] ),
    .QN(_13756_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01986_),
    .RN(net262),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.mscratch_q[15] ),
    .QN(_13755_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01987_),
    .RN(net265),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.mscratch_q[16] ),
    .QN(_13754_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01988_),
    .RN(net262),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.mscratch_q[17] ),
    .QN(_13753_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01989_),
    .RN(net265),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mscratch_q[18] ),
    .QN(_13752_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01990_),
    .RN(net262),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[19] ),
    .QN(_13751_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_01991_),
    .RN(net262),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[1] ),
    .QN(_13750_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01992_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[20] ),
    .QN(_13749_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01993_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.mscratch_q[21] ),
    .QN(_13748_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01994_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mscratch_q[22] ),
    .QN(_13747_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01995_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.mscratch_q[23] ),
    .QN(_13746_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01996_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mscratch_q[24] ),
    .QN(_13745_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01997_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mscratch_q[25] ),
    .QN(_13744_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01998_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[26] ),
    .QN(_13743_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01999_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[27] ),
    .QN(_13742_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02000_),
    .RN(net153),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mscratch_q[28] ),
    .QN(_13741_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02001_),
    .RN(net265),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[29] ),
    .QN(_13740_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02002_),
    .RN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mscratch_q[2] ),
    .QN(_13739_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02003_),
    .RN(net265),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mscratch_q[30] ),
    .QN(_13738_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02004_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[31] ),
    .QN(_13737_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02005_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.mscratch_q[3] ),
    .QN(_13736_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02006_),
    .RN(net262),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[4] ),
    .QN(_13735_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02007_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.mscratch_q[5] ),
    .QN(_13734_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02008_),
    .RN(net261),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mscratch_q[6] ),
    .QN(_13733_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02009_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.mscratch_q[7] ),
    .QN(_13732_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02010_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[8] ),
    .QN(_13731_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02011_),
    .RN(net265),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[9] ),
    .QN(_13730_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02012_),
    .RN(net262),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mstack_cause_q[0] ),
    .QN(_13729_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02013_),
    .RN(net262),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mstack_cause_q[1] ),
    .QN(_13728_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02014_),
    .RN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mstack_cause_q[2] ),
    .QN(_13727_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02015_),
    .RN(net265),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mstack_cause_q[3] ),
    .QN(_13726_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02016_),
    .RN(net265),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mstack_cause_q[4] ),
    .QN(_13725_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02017_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mstack_cause_q[5] ),
    .QN(_13724_));
 DFFR_X1 \cs_registers_i.u_mstack_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02018_),
    .RN(net262),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mstack_q[0] ),
    .QN(_13723_));
 DFFR_X1 \cs_registers_i.u_mstack_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02019_),
    .RN(net262),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mstack_q[1] ),
    .QN(_13722_));
 DFFS_X1 \cs_registers_i.u_mstack_csr.rdata_q[2]$_DFFE_PN1P_  (.D(_02020_),
    .SN(net262),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mstack_q[2] ),
    .QN(_13721_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02021_),
    .RN(net262),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mstack_epc_q[0] ),
    .QN(_13720_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02022_),
    .RN(net265),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.mstack_epc_q[10] ),
    .QN(_13719_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02023_),
    .RN(net264),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.mstack_epc_q[11] ),
    .QN(_13718_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02024_),
    .RN(net265),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.mstack_epc_q[12] ),
    .QN(_13717_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02025_),
    .RN(net265),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.mstack_epc_q[13] ),
    .QN(_13716_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02026_),
    .RN(net153),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mstack_epc_q[14] ),
    .QN(_13715_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02027_),
    .RN(net264),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.mstack_epc_q[15] ),
    .QN(_13714_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02028_),
    .RN(net153),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mstack_epc_q[16] ),
    .QN(_13713_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02029_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.mstack_epc_q[17] ),
    .QN(_13712_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02030_),
    .RN(net265),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.mstack_epc_q[18] ),
    .QN(_13711_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02031_),
    .RN(net265),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.mstack_epc_q[19] ),
    .QN(_13710_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02032_),
    .RN(net262),
    .CK(clknet_leaf_57_clk),
    .Q(\cs_registers_i.mstack_epc_q[1] ),
    .QN(_13709_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02033_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.mstack_epc_q[20] ),
    .QN(_13708_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02034_),
    .RN(net153),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mstack_epc_q[21] ),
    .QN(_13707_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02035_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.mstack_epc_q[22] ),
    .QN(_13706_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02036_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.mstack_epc_q[23] ),
    .QN(_13705_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02037_),
    .RN(net153),
    .CK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.mstack_epc_q[24] ),
    .QN(_13704_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02038_),
    .RN(net153),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mstack_epc_q[25] ),
    .QN(_13703_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02039_),
    .RN(net153),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.mstack_epc_q[26] ),
    .QN(_13702_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02040_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.mstack_epc_q[27] ),
    .QN(_13701_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02041_),
    .RN(net265),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.mstack_epc_q[28] ),
    .QN(_13700_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02042_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.mstack_epc_q[29] ),
    .QN(_13699_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02043_),
    .RN(net265),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mstack_epc_q[2] ),
    .QN(_13698_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02044_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[30] ),
    .QN(_13697_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02045_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.mstack_epc_q[31] ),
    .QN(_13696_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02046_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.mstack_epc_q[3] ),
    .QN(_13695_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02047_),
    .RN(net265),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mstack_epc_q[4] ),
    .QN(_13694_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02048_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.mstack_epc_q[5] ),
    .QN(_13693_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02049_),
    .RN(net265),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.mstack_epc_q[6] ),
    .QN(_13692_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02050_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.mstack_epc_q[7] ),
    .QN(_13691_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02051_),
    .RN(net264),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.mstack_epc_q[8] ),
    .QN(_13690_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02052_),
    .RN(net264),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.mstack_epc_q[9] ),
    .QN(_13689_));
 DFFR_X2 \cs_registers_i.u_mstatus_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02053_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.csr_mstatus_tw_o ),
    .QN(_13688_));
 DFFR_X1 \cs_registers_i.u_mstatus_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02054_),
    .RN(net262),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mstatus_q[1] ),
    .QN(_13687_));
 DFFR_X1 \cs_registers_i.u_mstatus_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02055_),
    .RN(net262),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.mstack_d[0] ),
    .QN(_13686_));
 DFFR_X2 \cs_registers_i.u_mstatus_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02056_),
    .RN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mstack_d[1] ),
    .QN(_13685_));
 DFFS_X2 \cs_registers_i.u_mstatus_csr.rdata_q[4]$_DFFE_PN1P_  (.D(_02057_),
    .SN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mstack_d[2] ),
    .QN(_13684_));
 DFFR_X2 \cs_registers_i.u_mstatus_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02058_),
    .RN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.csr_mstatus_mie_o ),
    .QN(_13683_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02059_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mtval_q[0] ),
    .QN(_13682_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02060_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.mtval_q[10] ),
    .QN(_13681_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02061_),
    .RN(net262),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[11] ),
    .QN(_13680_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02062_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[12] ),
    .QN(_13679_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02063_),
    .RN(net265),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mtval_q[13] ),
    .QN(_13678_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02064_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[14] ),
    .QN(_13677_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02065_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[15] ),
    .QN(_13676_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02066_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[16] ),
    .QN(_13675_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02067_),
    .RN(net262),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mtval_q[17] ),
    .QN(_13674_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02068_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[18] ),
    .QN(_13673_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02069_),
    .RN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mtval_q[19] ),
    .QN(_13672_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02070_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mtval_q[1] ),
    .QN(_13671_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02071_),
    .RN(net262),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.mtval_q[20] ),
    .QN(_13670_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02072_),
    .RN(net262),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mtval_q[21] ),
    .QN(_13669_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02073_),
    .RN(net265),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.mtval_q[22] ),
    .QN(_13668_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02074_),
    .RN(net262),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mtval_q[23] ),
    .QN(_13667_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02075_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.mtval_q[24] ),
    .QN(_13666_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02076_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mtval_q[25] ),
    .QN(_13665_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02077_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mtval_q[26] ),
    .QN(_13664_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02078_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mtval_q[27] ),
    .QN(_13663_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02079_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mtval_q[28] ),
    .QN(_13662_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02080_),
    .RN(net153),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mtval_q[29] ),
    .QN(_13661_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02081_),
    .RN(net262),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[2] ),
    .QN(_13660_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02082_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.mtval_q[30] ),
    .QN(_13659_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02083_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[31] ),
    .QN(_13658_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02084_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[3] ),
    .QN(_13657_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02085_),
    .RN(net262),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[4] ),
    .QN(_13656_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02086_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[5] ),
    .QN(_13655_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02087_),
    .RN(net262),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mtval_q[6] ),
    .QN(_13654_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02088_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[7] ),
    .QN(_13653_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02089_),
    .RN(net262),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[8] ),
    .QN(_13652_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02090_),
    .RN(net265),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mtval_q[9] ),
    .QN(_13651_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02091_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_mtvec_o[10] ),
    .QN(_01169_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02092_),
    .RN(net265),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.csr_mtvec_o[11] ),
    .QN(_00550_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02093_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_mtvec_o[12] ),
    .QN(_00549_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02094_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_mtvec_o[13] ),
    .QN(_01170_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02095_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_mtvec_o[14] ),
    .QN(_01171_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02096_),
    .RN(net265),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.csr_mtvec_o[15] ),
    .QN(_01172_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02097_),
    .RN(net153),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.csr_mtvec_o[16] ),
    .QN(_01173_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02098_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[17] ),
    .QN(_01174_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02099_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_mtvec_o[18] ),
    .QN(_01175_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02100_),
    .RN(net265),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_mtvec_o[19] ),
    .QN(_01176_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02101_),
    .RN(net153),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.csr_mtvec_o[20] ),
    .QN(_01177_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02102_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_mtvec_o[21] ),
    .QN(_01178_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02103_),
    .RN(net153),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[22] ),
    .QN(_01179_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02104_),
    .RN(net265),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_mtvec_o[23] ),
    .QN(_01180_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02105_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_mtvec_o[24] ),
    .QN(_01181_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02106_),
    .RN(net153),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.csr_mtvec_o[25] ),
    .QN(_01182_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02107_),
    .RN(net153),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[26] ),
    .QN(_01183_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02108_),
    .RN(net153),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[27] ),
    .QN(_00007_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02109_),
    .RN(net153),
    .CK(clknet_leaf_70_clk),
    .Q(\cs_registers_i.csr_mtvec_o[28] ),
    .QN(_00008_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02110_),
    .RN(net153),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.csr_mtvec_o[29] ),
    .QN(_00009_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02111_),
    .RN(net265),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[30] ),
    .QN(_00010_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02112_),
    .RN(net265),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[31] ),
    .QN(_00011_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02113_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[8] ),
    .QN(_01167_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02114_),
    .RN(net265),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[9] ),
    .QN(_01168_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_02115_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .QN(_13650_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_02116_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .QN(_15538_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_02117_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .QN(_15539_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_02118_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .QN(_00066_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_02119_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .QN(_00067_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_02120_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .QN(_01158_));
 DFFS_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .SN(net264),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .QN(_14051_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .RN(net264),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .QN(_00555_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .QN(_14052_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net264),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .QN(_14053_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .QN(_00178_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .QN(_13649_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_02121_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .QN(_00101_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_02122_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .QN(_00111_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_02123_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .QN(_00110_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_02124_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .QN(_00113_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_02125_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .QN(_00112_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_02126_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .QN(_00115_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_02127_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .QN(_00114_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_02128_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .QN(_00117_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_02129_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .QN(_00116_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_02130_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .QN(_00119_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_02131_),
    .RN(net263),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .QN(_00118_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_02132_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .QN(_00100_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_02133_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .QN(_00121_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_02134_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .QN(_00120_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_02135_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .QN(_00123_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_02136_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .QN(_00122_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_02137_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .QN(_00125_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_02138_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .QN(_00124_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_02139_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .QN(_00127_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_02140_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .QN(_00126_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_02141_),
    .RN(net263),
    .CK(clknet_leaf_13_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .QN(_00129_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_02142_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .QN(_00128_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_02143_),
    .RN(net263),
    .CK(clknet_leaf_11_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .QN(_00103_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_02144_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .QN(_00131_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_02145_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .QN(_00130_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_02146_),
    .RN(net263),
    .CK(clknet_leaf_12_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .QN(_00102_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_02147_),
    .RN(net263),
    .CK(clknet_leaf_11_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .QN(_00105_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_02148_),
    .RN(net263),
    .CK(clknet_leaf_11_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .QN(_00104_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_02149_),
    .RN(net263),
    .CK(clknet_leaf_11_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .QN(_00107_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_02150_),
    .RN(net263),
    .CK(clknet_leaf_11_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .QN(_00106_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_02151_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .QN(_00109_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_02152_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .QN(_00108_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_02153_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .QN(_00068_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_02154_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .QN(_00078_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_02155_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .QN(_00079_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_02156_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .QN(_00080_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_02157_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .QN(_00081_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_02158_),
    .RN(net264),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .QN(_00082_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_02159_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .QN(_00083_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_02160_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .QN(_00084_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_02161_),
    .RN(net264),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .QN(_00085_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_02162_),
    .RN(net264),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .QN(_00086_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_02163_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .QN(_00087_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_02164_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .QN(_00069_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_02165_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .QN(_00088_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_02166_),
    .RN(net264),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .QN(_00089_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_02167_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .QN(_00090_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_02168_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .QN(_00091_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_02169_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .QN(_00092_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_02170_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .QN(_00093_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_02171_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .QN(_00094_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_02172_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .QN(_00095_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_02173_),
    .RN(net264),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .QN(_00096_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_02174_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .QN(_00097_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_02175_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .QN(_00070_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_02176_),
    .RN(net264),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .QN(_00098_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_02177_),
    .RN(net264),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .QN(_00099_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_02178_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .QN(_00071_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_02179_),
    .RN(net264),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .QN(_00072_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_02180_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .QN(_00073_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_02181_),
    .RN(net264),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .QN(_00074_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_02182_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .QN(_00075_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_02183_),
    .RN(net264),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .QN(_00076_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_02184_),
    .RN(net264),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .QN(_00077_));
 DFFR_X1 \fetch_enable_q$_DFFE_PN0P_  (.D(_02185_),
    .RN(net261),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(fetch_enable_q),
    .QN(_13648_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[0]$_DFFE_PN0P_  (.D(_02186_),
    .RN(net259),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .QN(_13647_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[100]$_DFFE_PN0P_  (.D(_02187_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .QN(_00311_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[101]$_DFFE_PN0P_  (.D(_02188_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .QN(_00341_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[102]$_DFFE_PN0P_  (.D(_02189_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .QN(_00371_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[103]$_DFFE_PN0P_  (.D(_02190_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .QN(_00401_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[104]$_DFFE_PN0P_  (.D(_02191_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .QN(_00431_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[105]$_DFFE_PN0P_  (.D(_02192_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .QN(_00461_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[106]$_DFFE_PN0P_  (.D(_02193_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .QN(_00491_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[107]$_DFFE_PN0P_  (.D(_02194_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .QN(_00521_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[108]$_DFFE_PN0P_  (.D(_02195_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .QN(_00220_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[109]$_DFFE_PN0P_  (.D(_02196_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .QN(_00569_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[10]$_DFFE_PN0P_  (.D(_02197_),
    .RN(net256),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .QN(_13646_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[110]$_DFFE_PN0P_  (.D(_02198_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .QN(_00600_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[111]$_DFFE_PN0P_  (.D(_02199_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .QN(_00631_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[112]$_DFFE_PN0P_  (.D(_02200_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .QN(_00662_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[113]$_DFFE_PN0P_  (.D(_02201_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .QN(_00693_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[114]$_DFFE_PN0P_  (.D(_02202_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .QN(_00724_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[115]$_DFFE_PN0P_  (.D(_02203_),
    .RN(net260),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .QN(_00755_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[116]$_DFFE_PN0P_  (.D(_02204_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .QN(_00786_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[117]$_DFFE_PN0P_  (.D(_02205_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .QN(_00817_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[118]$_DFFE_PN0P_  (.D(_02206_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .QN(_00848_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[119]$_DFFE_PN0P_  (.D(_02207_),
    .RN(net258),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .QN(_00879_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[11]$_DFFE_PN0P_  (.D(_02208_),
    .RN(net263),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .QN(_13645_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[120]$_DFFE_PN0P_  (.D(_02209_),
    .RN(net258),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .QN(_00910_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[121]$_DFFE_PN0P_  (.D(_02210_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .QN(_00941_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[122]$_DFFE_PN0P_  (.D(_02211_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .QN(_00972_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[123]$_DFFE_PN0P_  (.D(_02212_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .QN(_01003_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[124]$_DFFE_PN0P_  (.D(_02213_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .QN(_01034_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[125]$_DFFE_PN0P_  (.D(_02214_),
    .RN(net258),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .QN(_01065_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[126]$_DFFE_PN0P_  (.D(_02215_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .QN(_01096_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[127]$_DFFE_PN0P_  (.D(_02216_),
    .RN(net259),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .QN(_01127_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[128]$_DFFE_PN0P_  (.D(_02217_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .QN(_00189_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[129]$_DFFE_PN0P_  (.D(_02218_),
    .RN(net259),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .QN(_00144_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[12]$_DFFE_PN0P_  (.D(_02219_),
    .RN(net256),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .QN(_13644_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[130]$_DFFE_PN0P_  (.D(_02220_),
    .RN(net259),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .QN(_00251_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[131]$_DFFE_PN0P_  (.D(_02221_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .QN(_00282_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[132]$_DFFE_PN0P_  (.D(_02222_),
    .RN(net263),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .QN(_00312_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[133]$_DFFE_PN0P_  (.D(_02223_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .QN(_00342_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[134]$_DFFE_PN0P_  (.D(_02224_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .QN(_00372_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[135]$_DFFE_PN0P_  (.D(_02225_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .QN(_00402_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[136]$_DFFE_PN0P_  (.D(_02226_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .QN(_00432_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[137]$_DFFE_PN0P_  (.D(_02227_),
    .RN(net263),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .QN(_00462_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[138]$_DFFE_PN0P_  (.D(_02228_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .QN(_00492_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[139]$_DFFE_PN0P_  (.D(_02229_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .QN(_00522_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[13]$_DFFE_PN0P_  (.D(_02230_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .QN(_13643_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[140]$_DFFE_PN0P_  (.D(_02231_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .QN(_00221_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[141]$_DFFE_PN0P_  (.D(_02232_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .QN(_00570_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[142]$_DFFE_PN0P_  (.D(_02233_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .QN(_00601_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[143]$_DFFE_PN0P_  (.D(_02234_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .QN(_00632_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[144]$_DFFE_PN0P_  (.D(_02235_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .QN(_00663_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[145]$_DFFE_PN0P_  (.D(_02236_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .QN(_00694_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[146]$_DFFE_PN0P_  (.D(_02237_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .QN(_00725_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[147]$_DFFE_PN0P_  (.D(_02238_),
    .RN(net259),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .QN(_00756_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[148]$_DFFE_PN0P_  (.D(_02239_),
    .RN(net258),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .QN(_00787_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[149]$_DFFE_PN0P_  (.D(_02240_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .QN(_00818_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[14]$_DFFE_PN0P_  (.D(_02241_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .QN(_13642_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[150]$_DFFE_PN0P_  (.D(_02242_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .QN(_00849_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[151]$_DFFE_PN0P_  (.D(_02243_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .QN(_00880_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[152]$_DFFE_PN0P_  (.D(_02244_),
    .RN(net258),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .QN(_00911_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[153]$_DFFE_PN0P_  (.D(_02245_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .QN(_00942_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[154]$_DFFE_PN0P_  (.D(_02246_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .QN(_00973_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[155]$_DFFE_PN0P_  (.D(_02247_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .QN(_01004_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[156]$_DFFE_PN0P_  (.D(_02248_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .QN(_01035_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[157]$_DFFE_PN0P_  (.D(_02249_),
    .RN(net258),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .QN(_01066_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[158]$_DFFE_PN0P_  (.D(_02250_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .QN(_01097_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[159]$_DFFE_PN0P_  (.D(_02251_),
    .RN(net259),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .QN(_01128_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[15]$_DFFE_PN0P_  (.D(_02252_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .QN(_13641_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[160]$_DFFE_PN0P_  (.D(_02253_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .QN(_00190_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[161]$_DFFE_PN0P_  (.D(_02254_),
    .RN(net259),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .QN(_00145_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[162]$_DFFE_PN0P_  (.D(_02255_),
    .RN(net259),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .QN(_00252_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[163]$_DFFE_PN0P_  (.D(_02256_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .QN(_00283_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[164]$_DFFE_PN0P_  (.D(_02257_),
    .RN(net263),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .QN(_00313_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[165]$_DFFE_PN0P_  (.D(_02258_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .QN(_00343_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[166]$_DFFE_PN0P_  (.D(_02259_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .QN(_00373_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[167]$_DFFE_PN0P_  (.D(_02260_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .QN(_00403_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[168]$_DFFE_PN0P_  (.D(_02261_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .QN(_00433_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[169]$_DFFE_PN0P_  (.D(_02262_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .QN(_00463_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[16]$_DFFE_PN0P_  (.D(_02263_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .QN(_13640_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[170]$_DFFE_PN0P_  (.D(_02264_),
    .RN(net256),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .QN(_00493_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[171]$_DFFE_PN0P_  (.D(_02265_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .QN(_00523_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[172]$_DFFE_PN0P_  (.D(_02266_),
    .RN(net260),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .QN(_00222_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[173]$_DFFE_PN0P_  (.D(_02267_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .QN(_00571_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[174]$_DFFE_PN0P_  (.D(_02268_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .QN(_00602_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[175]$_DFFE_PN0P_  (.D(_02269_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .QN(_00633_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[176]$_DFFE_PN0P_  (.D(_02270_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .QN(_00664_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[177]$_DFFE_PN0P_  (.D(_02271_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .QN(_00695_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[178]$_DFFE_PN0P_  (.D(_02272_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .QN(_00726_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[179]$_DFFE_PN0P_  (.D(_02273_),
    .RN(net258),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .QN(_00757_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[17]$_DFFE_PN0P_  (.D(_02274_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .QN(_13639_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[180]$_DFFE_PN0P_  (.D(_02275_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .QN(_00788_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[181]$_DFFE_PN0P_  (.D(_02276_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .QN(_00819_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[182]$_DFFE_PN0P_  (.D(_02277_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .QN(_00850_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[183]$_DFFE_PN0P_  (.D(_02278_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .QN(_00881_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[184]$_DFFE_PN0P_  (.D(_02279_),
    .RN(net260),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .QN(_00912_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[185]$_DFFE_PN0P_  (.D(_02280_),
    .RN(net260),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .QN(_00943_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[186]$_DFFE_PN0P_  (.D(_02281_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .QN(_00974_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[187]$_DFFE_PN0P_  (.D(_02282_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .QN(_01005_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[188]$_DFFE_PN0P_  (.D(_02283_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .QN(_01036_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[189]$_DFFE_PN0P_  (.D(_02284_),
    .RN(net258),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .QN(_01067_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[18]$_DFFE_PN0P_  (.D(_02285_),
    .RN(net257),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .QN(_13638_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[190]$_DFFE_PN0P_  (.D(_02286_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .QN(_01098_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[191]$_DFFE_PN0P_  (.D(_02287_),
    .RN(net260),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .QN(_01129_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[192]$_DFFE_PN0P_  (.D(_02288_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .QN(_00191_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[193]$_DFFE_PN0P_  (.D(_02289_),
    .RN(net259),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .QN(_00146_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[194]$_DFFE_PN0P_  (.D(_02290_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .QN(_00253_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[195]$_DFFE_PN0P_  (.D(_02291_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .QN(_00284_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[196]$_DFFE_PN0P_  (.D(_02292_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .QN(_00314_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[197]$_DFFE_PN0P_  (.D(_02293_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .QN(_00344_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[198]$_DFFE_PN0P_  (.D(_02294_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .QN(_00374_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[199]$_DFFE_PN0P_  (.D(_02295_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .QN(_00404_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[19]$_DFFE_PN0P_  (.D(_02296_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .QN(_13637_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[1]$_DFFE_PN0P_  (.D(_02297_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .QN(_13636_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[200]$_DFFE_PN0P_  (.D(_02298_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .QN(_00434_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[201]$_DFFE_PN0P_  (.D(_02299_),
    .RN(net263),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .QN(_00464_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[202]$_DFFE_PN0P_  (.D(_02300_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .QN(_00494_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[203]$_DFFE_PN0P_  (.D(_02301_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .QN(_00524_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[204]$_DFFE_PN0P_  (.D(_02302_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .QN(_00223_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[205]$_DFFE_PN0P_  (.D(_02303_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .QN(_00572_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[206]$_DFFE_PN0P_  (.D(_02304_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .QN(_00603_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[207]$_DFFE_PN0P_  (.D(_02305_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .QN(_00634_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[208]$_DFFE_PN0P_  (.D(_02306_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .QN(_00665_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[209]$_DFFE_PN0P_  (.D(_02307_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .QN(_00696_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[20]$_DFFE_PN0P_  (.D(_02308_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .QN(_13635_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[210]$_DFFE_PN0P_  (.D(_02309_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .QN(_00727_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[211]$_DFFE_PN0P_  (.D(_02310_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .QN(_00758_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[212]$_DFFE_PN0P_  (.D(_02311_),
    .RN(net258),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .QN(_00789_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[213]$_DFFE_PN0P_  (.D(_02312_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .QN(_00820_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[214]$_DFFE_PN0P_  (.D(_02313_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .QN(_00851_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[215]$_DFFE_PN0P_  (.D(_02314_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .QN(_00882_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[216]$_DFFE_PN0P_  (.D(_02315_),
    .RN(net258),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .QN(_00913_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[217]$_DFFE_PN0P_  (.D(_02316_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .QN(_00944_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[218]$_DFFE_PN0P_  (.D(_02317_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .QN(_00975_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[219]$_DFFE_PN0P_  (.D(_02318_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .QN(_01006_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[21]$_DFFE_PN0P_  (.D(_02319_),
    .RN(net260),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .QN(_13634_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[220]$_DFFE_PN0P_  (.D(_02320_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .QN(_01037_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[221]$_DFFE_PN0P_  (.D(_02321_),
    .RN(net258),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .QN(_01068_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[222]$_DFFE_PN0P_  (.D(_02322_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .QN(_01099_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[223]$_DFFE_PN0P_  (.D(_02323_),
    .RN(net259),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .QN(_01130_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[224]$_DFFE_PN0P_  (.D(_02324_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .QN(_00192_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[225]$_DFFE_PN0P_  (.D(_02325_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .QN(_00147_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[226]$_DFFE_PN0P_  (.D(_02326_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .QN(_00254_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[227]$_DFFE_PN0P_  (.D(_02327_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .QN(_00285_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[228]$_DFFE_PN0P_  (.D(_02328_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .QN(_00315_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[229]$_DFFE_PN0P_  (.D(_02329_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .QN(_00345_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[22]$_DFFE_PN0P_  (.D(_02330_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .QN(_13633_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[230]$_DFFE_PN0P_  (.D(_02331_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .QN(_00375_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[231]$_DFFE_PN0P_  (.D(_02332_),
    .RN(net263),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .QN(_00405_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[232]$_DFFE_PN0P_  (.D(_02333_),
    .RN(net259),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .QN(_00435_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[233]$_DFFE_PN0P_  (.D(_02334_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .QN(_00465_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[234]$_DFFE_PN0P_  (.D(_02335_),
    .RN(net256),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .QN(_00495_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[235]$_DFFE_PN0P_  (.D(_02336_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .QN(_00525_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[236]$_DFFE_PN0P_  (.D(_02337_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .QN(_00224_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[237]$_DFFE_PN0P_  (.D(_02338_),
    .RN(net256),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .QN(_00573_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[238]$_DFFE_PN0P_  (.D(_02339_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .QN(_00604_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[239]$_DFFE_PN0P_  (.D(_02340_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .QN(_00635_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[23]$_DFFE_PN0P_  (.D(_02341_),
    .RN(net258),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .QN(_13632_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[240]$_DFFE_PN0P_  (.D(_02342_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .QN(_00666_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[241]$_DFFE_PN0P_  (.D(_02343_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .QN(_00697_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[242]$_DFFE_PN0P_  (.D(_02344_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .QN(_00728_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[243]$_DFFE_PN0P_  (.D(_02345_),
    .RN(net260),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .QN(_00759_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[244]$_DFFE_PN0P_  (.D(_02346_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .QN(_00790_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[245]$_DFFE_PN0P_  (.D(_02347_),
    .RN(net260),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .QN(_00821_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[246]$_DFFE_PN0P_  (.D(_02348_),
    .RN(net258),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .QN(_00852_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[247]$_DFFE_PN0P_  (.D(_02349_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .QN(_00883_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[248]$_DFFE_PN0P_  (.D(_02350_),
    .RN(net260),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .QN(_00914_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[249]$_DFFE_PN0P_  (.D(_02351_),
    .RN(net260),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .QN(_00945_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[24]$_DFFE_PN0P_  (.D(_02352_),
    .RN(net260),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .QN(_13631_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[250]$_DFFE_PN0P_  (.D(_02353_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .QN(_00976_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[251]$_DFFE_PN0P_  (.D(_02354_),
    .RN(net258),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .QN(_01007_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[252]$_DFFE_PN0P_  (.D(_02355_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .QN(_01038_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[253]$_DFFE_PN0P_  (.D(_02356_),
    .RN(net260),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .QN(_01069_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[254]$_DFFE_PN0P_  (.D(_02357_),
    .RN(net260),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .QN(_01100_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[255]$_DFFE_PN0P_  (.D(_02358_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .QN(_01131_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[256]$_DFFE_PN0P_  (.D(_02359_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .QN(_00193_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[257]$_DFFE_PN0P_  (.D(_02360_),
    .RN(net259),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .QN(_00148_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[258]$_DFFE_PN0P_  (.D(_02361_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .QN(_00255_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[259]$_DFFE_PN0P_  (.D(_02362_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .QN(_00286_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[25]$_DFFE_PN0P_  (.D(_02363_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .QN(_13630_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[260]$_DFFE_PN0P_  (.D(_02364_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .QN(_00316_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[261]$_DFFE_PN0P_  (.D(_02365_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .QN(_00346_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[262]$_DFFE_PN0P_  (.D(_02366_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .QN(_00376_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[263]$_DFFE_PN0P_  (.D(_02367_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .QN(_00406_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[264]$_DFFE_PN0P_  (.D(_02368_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .QN(_00436_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[265]$_DFFE_PN0P_  (.D(_02369_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .QN(_00466_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[266]$_DFFE_PN0P_  (.D(_02370_),
    .RN(net256),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .QN(_00496_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[267]$_DFFE_PN0P_  (.D(_02371_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .QN(_00526_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[268]$_DFFE_PN0P_  (.D(_02372_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .QN(_00225_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[269]$_DFFE_PN0P_  (.D(_02373_),
    .RN(net256),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .QN(_00574_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[26]$_DFFE_PN0P_  (.D(_02374_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .QN(_13629_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[270]$_DFFE_PN0P_  (.D(_02375_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .QN(_00605_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[271]$_DFFE_PN0P_  (.D(_02376_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .QN(_00636_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[272]$_DFFE_PN0P_  (.D(_02377_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .QN(_00667_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[273]$_DFFE_PN0P_  (.D(_02378_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .QN(_00698_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[274]$_DFFE_PN0P_  (.D(_02379_),
    .RN(net256),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .QN(_00729_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[275]$_DFFE_PN0P_  (.D(_02380_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .QN(_00760_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[276]$_DFFE_PN0P_  (.D(_02381_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .QN(_00791_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[277]$_DFFE_PN0P_  (.D(_02382_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .QN(_00822_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[278]$_DFFE_PN0P_  (.D(_02383_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .QN(_00853_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[279]$_DFFE_PN0P_  (.D(_02384_),
    .RN(net258),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .QN(_00884_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[27]$_DFFE_PN0P_  (.D(_02385_),
    .RN(net260),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .QN(_13628_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[280]$_DFFE_PN0P_  (.D(_02386_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .QN(_00915_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[281]$_DFFE_PN0P_  (.D(_02387_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .QN(_00946_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[282]$_DFFE_PN0P_  (.D(_02388_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .QN(_00977_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[283]$_DFFE_PN0P_  (.D(_02389_),
    .RN(net258),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .QN(_01008_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[284]$_DFFE_PN0P_  (.D(_02390_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .QN(_01039_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[285]$_DFFE_PN0P_  (.D(_02391_),
    .RN(net258),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .QN(_01070_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[286]$_DFFE_PN0P_  (.D(_02392_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .QN(_01101_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[287]$_DFFE_PN0P_  (.D(_02393_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .QN(_01132_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[288]$_DFFE_PN0P_  (.D(_02394_),
    .RN(net259),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .QN(_00194_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[289]$_DFFE_PN0P_  (.D(_02395_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .QN(_00149_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[28]$_DFFE_PN0P_  (.D(_02396_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .QN(_13627_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[290]$_DFFE_PN0P_  (.D(_02397_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .QN(_00256_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[291]$_DFFE_PN0P_  (.D(_02398_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .QN(_00287_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[292]$_DFFE_PN0P_  (.D(_02399_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .QN(_00317_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[293]$_DFFE_PN0P_  (.D(_02400_),
    .RN(net259),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .QN(_00347_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[294]$_DFFE_PN0P_  (.D(_02401_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .QN(_00377_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[295]$_DFFE_PN0P_  (.D(_02402_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .QN(_00407_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[296]$_DFFE_PN0P_  (.D(_02403_),
    .RN(net259),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .QN(_00437_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[297]$_DFFE_PN0P_  (.D(_02404_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .QN(_00467_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[298]$_DFFE_PN0P_  (.D(_02405_),
    .RN(net256),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .QN(_00497_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[299]$_DFFE_PN0P_  (.D(_02406_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .QN(_00527_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[29]$_DFFE_PN0P_  (.D(_02407_),
    .RN(net259),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .QN(_13626_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[2]$_DFFE_PN0P_  (.D(_02408_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .QN(_13625_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[300]$_DFFE_PN0P_  (.D(_02409_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .QN(_00226_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[301]$_DFFE_PN0P_  (.D(_02410_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .QN(_00575_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[302]$_DFFE_PN0P_  (.D(_02411_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .QN(_00606_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[303]$_DFFE_PN0P_  (.D(_02412_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .QN(_00637_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[304]$_DFFE_PN0P_  (.D(_02413_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .QN(_00668_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[305]$_DFFE_PN0P_  (.D(_02414_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .QN(_00699_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[306]$_DFFE_PN0P_  (.D(_02415_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .QN(_00730_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[307]$_DFFE_PN0P_  (.D(_02416_),
    .RN(net260),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .QN(_00761_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[308]$_DFFE_PN0P_  (.D(_02417_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .QN(_00792_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[309]$_DFFE_PN0P_  (.D(_02418_),
    .RN(net260),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .QN(_00823_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[30]$_DFFE_PN0P_  (.D(_02419_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .QN(_13624_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[310]$_DFFE_PN0P_  (.D(_02420_),
    .RN(net258),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .QN(_00854_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[311]$_DFFE_PN0P_  (.D(_02421_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .QN(_00885_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[312]$_DFFE_PN0P_  (.D(_02422_),
    .RN(net260),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .QN(_00916_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[313]$_DFFE_PN0P_  (.D(_02423_),
    .RN(net260),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .QN(_00947_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[314]$_DFFE_PN0P_  (.D(_02424_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .QN(_00978_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[315]$_DFFE_PN0P_  (.D(_02425_),
    .RN(net258),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .QN(_01009_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[316]$_DFFE_PN0P_  (.D(_02426_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .QN(_01040_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[317]$_DFFE_PN0P_  (.D(_02427_),
    .RN(net260),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .QN(_01071_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[318]$_DFFE_PN0P_  (.D(_02428_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .QN(_01102_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[319]$_DFFE_PN0P_  (.D(_02429_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .QN(_01133_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[31]$_DFFE_PN0P_  (.D(_02430_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .QN(_13623_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[320]$_DFFE_PN0P_  (.D(_02431_),
    .RN(net259),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .QN(_00195_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[321]$_DFFE_PN0P_  (.D(_02432_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .QN(_00150_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[322]$_DFFE_PN0P_  (.D(_02433_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .QN(_00257_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[323]$_DFFE_PN0P_  (.D(_02434_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .QN(_00288_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[324]$_DFFE_PN0P_  (.D(_02435_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .QN(_00318_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[325]$_DFFE_PN0P_  (.D(_02436_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .QN(_00348_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[326]$_DFFE_PN0P_  (.D(_02437_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .QN(_00378_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[327]$_DFFE_PN0P_  (.D(_02438_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .QN(_00408_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[328]$_DFFE_PN0P_  (.D(_02439_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .QN(_00438_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[329]$_DFFE_PN0P_  (.D(_02440_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .QN(_00468_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[32]$_DFFE_PN0P_  (.D(_02441_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .QN(_00186_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[330]$_DFFE_PN0P_  (.D(_02442_),
    .RN(net256),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .QN(_00498_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[331]$_DFFE_PN0P_  (.D(_02443_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .QN(_00528_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[332]$_DFFE_PN0P_  (.D(_02444_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .QN(_00227_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[333]$_DFFE_PN0P_  (.D(_02445_),
    .RN(net256),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .QN(_00576_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[334]$_DFFE_PN0P_  (.D(_02446_),
    .RN(net257),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .QN(_00607_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[335]$_DFFE_PN0P_  (.D(_02447_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .QN(_00638_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[336]$_DFFE_PN0P_  (.D(_02448_),
    .RN(net257),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .QN(_00669_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[337]$_DFFE_PN0P_  (.D(_02449_),
    .RN(net257),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .QN(_00700_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[338]$_DFFE_PN0P_  (.D(_02450_),
    .RN(net256),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .QN(_00731_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[339]$_DFFE_PN0P_  (.D(_02451_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .QN(_00762_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[33]$_DFFE_PN0P_  (.D(_02452_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .QN(_00141_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[340]$_DFFE_PN0P_  (.D(_02453_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .QN(_00793_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[341]$_DFFE_PN0P_  (.D(_02454_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .QN(_00824_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[342]$_DFFE_PN0P_  (.D(_02455_),
    .RN(net258),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .QN(_00855_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[343]$_DFFE_PN0P_  (.D(_02456_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .QN(_00886_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[344]$_DFFE_PN0P_  (.D(_02457_),
    .RN(net260),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .QN(_00917_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[345]$_DFFE_PN0P_  (.D(_02458_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .QN(_00948_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[346]$_DFFE_PN0P_  (.D(_02459_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .QN(_00979_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[347]$_DFFE_PN0P_  (.D(_02460_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .QN(_01010_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[348]$_DFFE_PN0P_  (.D(_02461_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .QN(_01041_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[349]$_DFFE_PN0P_  (.D(_02462_),
    .RN(net260),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .QN(_01072_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[34]$_DFFE_PN0P_  (.D(_02463_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .QN(_00248_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[350]$_DFFE_PN0P_  (.D(_02464_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .QN(_01103_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[351]$_DFFE_PN0P_  (.D(_02465_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .QN(_01134_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[352]$_DFFE_PN0P_  (.D(_02466_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .QN(_00196_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[353]$_DFFE_PN0P_  (.D(_02467_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .QN(_00151_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[354]$_DFFE_PN0P_  (.D(_02468_),
    .RN(net256),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .QN(_00258_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[355]$_DFFE_PN0P_  (.D(_02469_),
    .RN(net256),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .QN(_00289_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[356]$_DFFE_PN0P_  (.D(_02470_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .QN(_00319_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[357]$_DFFE_PN0P_  (.D(_02471_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .QN(_00349_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[358]$_DFFE_PN0P_  (.D(_02472_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .QN(_00379_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[359]$_DFFE_PN0P_  (.D(_02473_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .QN(_00409_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[35]$_DFFE_PN0P_  (.D(_02474_),
    .RN(net259),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .QN(_00279_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[360]$_DFFE_PN0P_  (.D(_02475_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .QN(_00439_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[361]$_DFFE_PN0P_  (.D(_02476_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .QN(_00469_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[362]$_DFFE_PN0P_  (.D(_02477_),
    .RN(net256),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .QN(_00499_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[363]$_DFFE_PN0P_  (.D(_02478_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .QN(_00529_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[364]$_DFFE_PN0P_  (.D(_02479_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .QN(_00228_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[365]$_DFFE_PN0P_  (.D(_02480_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .QN(_00577_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[366]$_DFFE_PN0P_  (.D(_02481_),
    .RN(net257),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .QN(_00608_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[367]$_DFFE_PN0P_  (.D(_02482_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .QN(_00639_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[368]$_DFFE_PN0P_  (.D(_02483_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .QN(_00670_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[369]$_DFFE_PN0P_  (.D(_02484_),
    .RN(net260),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .QN(_00701_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[36]$_DFFE_PN0P_  (.D(_02485_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .QN(_00309_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[370]$_DFFE_PN0P_  (.D(_02486_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .QN(_00732_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[371]$_DFFE_PN0P_  (.D(_02487_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .QN(_00763_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[372]$_DFFE_PN0P_  (.D(_02488_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .QN(_00794_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[373]$_DFFE_PN0P_  (.D(_02489_),
    .RN(net258),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .QN(_00825_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[374]$_DFFE_PN0P_  (.D(_02490_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .QN(_00856_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[375]$_DFFE_PN0P_  (.D(_02491_),
    .RN(net255),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .QN(_00887_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[376]$_DFFE_PN0P_  (.D(_02492_),
    .RN(net258),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .QN(_00918_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[377]$_DFFE_PN0P_  (.D(_02493_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .QN(_00949_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[378]$_DFFE_PN0P_  (.D(_02494_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .QN(_00980_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[379]$_DFFE_PN0P_  (.D(_02495_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .QN(_01011_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[37]$_DFFE_PN0P_  (.D(_02496_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .QN(_00339_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[380]$_DFFE_PN0P_  (.D(_02497_),
    .RN(net258),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .QN(_01042_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[381]$_DFFE_PN0P_  (.D(_02498_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .QN(_01073_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[382]$_DFFE_PN0P_  (.D(_02499_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .QN(_01104_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[383]$_DFFE_PN0P_  (.D(_02500_),
    .RN(net259),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .QN(_01135_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[384]$_DFFE_PN0P_  (.D(_02501_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .QN(_00197_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[385]$_DFFE_PN0P_  (.D(_02502_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .QN(_00152_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[386]$_DFFE_PN0P_  (.D(_02503_),
    .RN(net256),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .QN(_00259_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[387]$_DFFE_PN0P_  (.D(_02504_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .QN(_00290_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[388]$_DFFE_PN0P_  (.D(_02505_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .QN(_00320_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[389]$_DFFE_PN0P_  (.D(_02506_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .QN(_00350_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[38]$_DFFE_PN0P_  (.D(_02507_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .QN(_00369_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[390]$_DFFE_PN0P_  (.D(_02508_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .QN(_00380_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[391]$_DFFE_PN0P_  (.D(_02509_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .QN(_00410_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[392]$_DFFE_PN0P_  (.D(_02510_),
    .RN(net259),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .QN(_00440_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[393]$_DFFE_PN0P_  (.D(_02511_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .QN(_00470_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[394]$_DFFE_PN0P_  (.D(_02512_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .QN(_00500_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[395]$_DFFE_PN0P_  (.D(_02513_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .QN(_00530_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[396]$_DFFE_PN0P_  (.D(_02514_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .QN(_00229_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[397]$_DFFE_PN0P_  (.D(_02515_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .QN(_00578_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[398]$_DFFE_PN0P_  (.D(_02516_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .QN(_00609_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[399]$_DFFE_PN0P_  (.D(_02517_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .QN(_00640_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[39]$_DFFE_PN0P_  (.D(_02518_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .QN(_00399_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[3]$_DFFE_PN0P_  (.D(_02519_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .QN(_13622_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[400]$_DFFE_PN0P_  (.D(_02520_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .QN(_00671_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[401]$_DFFE_PN0P_  (.D(_02521_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .QN(_00702_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[402]$_DFFE_PN0P_  (.D(_02522_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .QN(_00733_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[403]$_DFFE_PN0P_  (.D(_02523_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .QN(_00764_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[404]$_DFFE_PN0P_  (.D(_02524_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .QN(_00795_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[405]$_DFFE_PN0P_  (.D(_02525_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .QN(_00826_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[406]$_DFFE_PN0P_  (.D(_02526_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .QN(_00857_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[407]$_DFFE_PN0P_  (.D(_02527_),
    .RN(net255),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .QN(_00888_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[408]$_DFFE_PN0P_  (.D(_02528_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .QN(_00919_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[409]$_DFFE_PN0P_  (.D(_02529_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .QN(_00950_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[40]$_DFFE_PN0P_  (.D(_02530_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .QN(_00429_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[410]$_DFFE_PN0P_  (.D(_02531_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .QN(_00981_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[411]$_DFFE_PN0P_  (.D(_02532_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .QN(_01012_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[412]$_DFFE_PN0P_  (.D(_02533_),
    .RN(net258),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .QN(_01043_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[413]$_DFFE_PN0P_  (.D(_02534_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .QN(_01074_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[414]$_DFFE_PN0P_  (.D(_02535_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .QN(_01105_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[415]$_DFFE_PN0P_  (.D(_02536_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .QN(_01136_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[416]$_DFFE_PN0P_  (.D(_02537_),
    .RN(net259),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .QN(_00198_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[417]$_DFFE_PN0P_  (.D(_02538_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .QN(_00153_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[418]$_DFFE_PN0P_  (.D(_02539_),
    .RN(net256),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .QN(_00260_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[419]$_DFFE_PN0P_  (.D(_02540_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .QN(_00291_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[41]$_DFFE_PN0P_  (.D(_02541_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .QN(_00459_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[420]$_DFFE_PN0P_  (.D(_02542_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .QN(_00321_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[421]$_DFFE_PN0P_  (.D(_02543_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .QN(_00351_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[422]$_DFFE_PN0P_  (.D(_02544_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .QN(_00381_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[423]$_DFFE_PN0P_  (.D(_02545_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .QN(_00411_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[424]$_DFFE_PN0P_  (.D(_02546_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .QN(_00441_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[425]$_DFFE_PN0P_  (.D(_02547_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .QN(_00471_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[426]$_DFFE_PN0P_  (.D(_02548_),
    .RN(net256),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .QN(_00501_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[427]$_DFFE_PN0P_  (.D(_02549_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .QN(_00531_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[428]$_DFFE_PN0P_  (.D(_02550_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .QN(_00230_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[429]$_DFFE_PN0P_  (.D(_02551_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .QN(_00579_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[42]$_DFFE_PN0P_  (.D(_02552_),
    .RN(net256),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .QN(_00489_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[430]$_DFFE_PN0P_  (.D(_02553_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .QN(_00610_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[431]$_DFFE_PN0P_  (.D(_02554_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .QN(_00641_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[432]$_DFFE_PN0P_  (.D(_02555_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .QN(_00672_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[433]$_DFFE_PN0P_  (.D(_02556_),
    .RN(net260),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .QN(_00703_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[434]$_DFFE_PN0P_  (.D(_02557_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .QN(_00734_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[435]$_DFFE_PN0P_  (.D(_02558_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .QN(_00765_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[436]$_DFFE_PN0P_  (.D(_02559_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .QN(_00796_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[437]$_DFFE_PN0P_  (.D(_02560_),
    .RN(net258),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .QN(_00827_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[438]$_DFFE_PN0P_  (.D(_02561_),
    .RN(net258),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .QN(_00858_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[439]$_DFFE_PN0P_  (.D(_02562_),
    .RN(net258),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .QN(_00889_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[43]$_DFFE_PN0P_  (.D(_02563_),
    .RN(net263),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .QN(_00519_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[440]$_DFFE_PN0P_  (.D(_02564_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .QN(_00920_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[441]$_DFFE_PN0P_  (.D(_02565_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .QN(_00951_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[442]$_DFFE_PN0P_  (.D(_02566_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .QN(_00982_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[443]$_DFFE_PN0P_  (.D(_02567_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .QN(_01013_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[444]$_DFFE_PN0P_  (.D(_02568_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .QN(_01044_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[445]$_DFFE_PN0P_  (.D(_02569_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .QN(_01075_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[446]$_DFFE_PN0P_  (.D(_02570_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .QN(_01106_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[447]$_DFFE_PN0P_  (.D(_02571_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .QN(_01137_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[448]$_DFFE_PN0P_  (.D(_02572_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .QN(_00199_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[449]$_DFFE_PN0P_  (.D(_02573_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .QN(_00154_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[44]$_DFFE_PN0P_  (.D(_02574_),
    .RN(net256),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .QN(_00218_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[450]$_DFFE_PN0P_  (.D(_02575_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .QN(_00261_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[451]$_DFFE_PN0P_  (.D(_02576_),
    .RN(net256),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .QN(_00292_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[452]$_DFFE_PN0P_  (.D(_02577_),
    .RN(net263),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .QN(_00322_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[453]$_DFFE_PN0P_  (.D(_02578_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .QN(_00352_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[454]$_DFFE_PN0P_  (.D(_02579_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .QN(_00382_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[455]$_DFFE_PN0P_  (.D(_02580_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .QN(_00412_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[456]$_DFFE_PN0P_  (.D(_02581_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .QN(_00442_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[457]$_DFFE_PN0P_  (.D(_02582_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .QN(_00472_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[458]$_DFFE_PN0P_  (.D(_02583_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .QN(_00502_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[459]$_DFFE_PN0P_  (.D(_02584_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .QN(_00532_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[45]$_DFFE_PN0P_  (.D(_02585_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .QN(_00567_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[460]$_DFFE_PN0P_  (.D(_02586_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .QN(_00231_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[461]$_DFFE_PN0P_  (.D(_02587_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .QN(_00580_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[462]$_DFFE_PN0P_  (.D(_02588_),
    .RN(net257),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .QN(_00611_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[463]$_DFFE_PN0P_  (.D(_02589_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .QN(_00642_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[464]$_DFFE_PN0P_  (.D(_02590_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .QN(_00673_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[465]$_DFFE_PN0P_  (.D(_02591_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .QN(_00704_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[466]$_DFFE_PN0P_  (.D(_02592_),
    .RN(net257),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .QN(_00735_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[467]$_DFFE_PN0P_  (.D(_02593_),
    .RN(net260),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .QN(_00766_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[468]$_DFFE_PN0P_  (.D(_02594_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .QN(_00797_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[469]$_DFFE_PN0P_  (.D(_02595_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .QN(_00828_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[46]$_DFFE_PN0P_  (.D(_02596_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .QN(_00598_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[470]$_DFFE_PN0P_  (.D(_02597_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .QN(_00859_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[471]$_DFFE_PN0P_  (.D(_02598_),
    .RN(net258),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .QN(_00890_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[472]$_DFFE_PN0P_  (.D(_02599_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .QN(_00921_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[473]$_DFFE_PN0P_  (.D(_02600_),
    .RN(net260),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .QN(_00952_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[474]$_DFFE_PN0P_  (.D(_02601_),
    .RN(net255),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .QN(_00983_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[475]$_DFFE_PN0P_  (.D(_02602_),
    .RN(net258),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .QN(_01014_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[476]$_DFFE_PN0P_  (.D(_02603_),
    .RN(net258),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .QN(_01045_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[477]$_DFFE_PN0P_  (.D(_02604_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .QN(_01076_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[478]$_DFFE_PN0P_  (.D(_02605_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .QN(_01107_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[479]$_DFFE_PN0P_  (.D(_02606_),
    .RN(net259),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .QN(_01138_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[47]$_DFFE_PN0P_  (.D(_02607_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .QN(_00629_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[480]$_DFFE_PN0P_  (.D(_02608_),
    .RN(net259),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .QN(_00200_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[481]$_DFFE_PN0P_  (.D(_02609_),
    .RN(net259),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .QN(_00155_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[482]$_DFFE_PN0P_  (.D(_02610_),
    .RN(net259),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .QN(_00262_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[483]$_DFFE_PN0P_  (.D(_02611_),
    .RN(net259),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .QN(_00293_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[484]$_DFFE_PN0P_  (.D(_02612_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .QN(_00323_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[485]$_DFFE_PN0P_  (.D(_02613_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .QN(_00353_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[486]$_DFFE_PN0P_  (.D(_02614_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .QN(_00383_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[487]$_DFFE_PN0P_  (.D(_02615_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .QN(_00413_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[488]$_DFFE_PN0P_  (.D(_02616_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .QN(_00443_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[489]$_DFFE_PN0P_  (.D(_02617_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .QN(_00473_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[48]$_DFFE_PN0P_  (.D(_02618_),
    .RN(net257),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .QN(_00660_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[490]$_DFFE_PN0P_  (.D(_02619_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .QN(_00503_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[491]$_DFFE_PN0P_  (.D(_02620_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .QN(_00533_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[492]$_DFFE_PN0P_  (.D(_02621_),
    .RN(net259),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .QN(_00232_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[493]$_DFFE_PN0P_  (.D(_02622_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .QN(_00581_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[494]$_DFFE_PN0P_  (.D(_02623_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .QN(_00612_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[495]$_DFFE_PN0P_  (.D(_02624_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .QN(_00643_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[496]$_DFFE_PN0P_  (.D(_02625_),
    .RN(net257),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .QN(_00674_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[497]$_DFFE_PN0P_  (.D(_02626_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .QN(_00705_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[498]$_DFFE_PN0P_  (.D(_02627_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .QN(_00736_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[499]$_DFFE_PN0P_  (.D(_02628_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .QN(_00767_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[49]$_DFFE_PN0P_  (.D(_02629_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .QN(_00691_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[4]$_DFFE_PN0P_  (.D(_02630_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .QN(_13621_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[500]$_DFFE_PN0P_  (.D(_02631_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .QN(_00798_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[501]$_DFFE_PN0P_  (.D(_02632_),
    .RN(net258),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .QN(_00829_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[502]$_DFFE_PN0P_  (.D(_02633_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .QN(_00860_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[503]$_DFFE_PN0P_  (.D(_02634_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .QN(_00891_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[504]$_DFFE_PN0P_  (.D(_02635_),
    .RN(net260),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .QN(_00922_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[505]$_DFFE_PN0P_  (.D(_02636_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .QN(_00953_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[506]$_DFFE_PN0P_  (.D(_02637_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .QN(_00984_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[507]$_DFFE_PN0P_  (.D(_02638_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .QN(_01015_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[508]$_DFFE_PN0P_  (.D(_02639_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .QN(_01046_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[509]$_DFFE_PN0P_  (.D(_02640_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .QN(_01077_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[50]$_DFFE_PN0P_  (.D(_02641_),
    .RN(net256),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .QN(_00722_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[510]$_DFFE_PN0P_  (.D(_02642_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .QN(_01108_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[511]$_DFFE_PN0P_  (.D(_02643_),
    .RN(net260),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .QN(_01139_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[512]$_DFFE_PN0P_  (.D(_02644_),
    .RN(net256),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .QN(_00201_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[513]$_DFFE_PN0P_  (.D(_02645_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .QN(_00156_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[514]$_DFFE_PN0P_  (.D(_02646_),
    .RN(net259),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .QN(_00263_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[515]$_DFFE_PN0P_  (.D(_02647_),
    .RN(net259),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .QN(_00294_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[516]$_DFFE_PN0P_  (.D(_02648_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .QN(_00324_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[517]$_DFFE_PN0P_  (.D(_02649_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .QN(_00354_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[518]$_DFFE_PN0P_  (.D(_02650_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .QN(_00384_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[519]$_DFFE_PN0P_  (.D(_02651_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .QN(_00414_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[51]$_DFFE_PN0P_  (.D(_02652_),
    .RN(net260),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .QN(_00753_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[520]$_DFFE_PN0P_  (.D(_02653_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .QN(_00444_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[521]$_DFFE_PN0P_  (.D(_02654_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .QN(_00474_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[522]$_DFFE_PN0P_  (.D(_02655_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .QN(_00504_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[523]$_DFFE_PN0P_  (.D(_02656_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .QN(_00534_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[524]$_DFFE_PN0P_  (.D(_02657_),
    .RN(net259),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .QN(_00233_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[525]$_DFFE_PN0P_  (.D(_02658_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .QN(_00582_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[526]$_DFFE_PN0P_  (.D(_02659_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .QN(_00613_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[527]$_DFFE_PN0P_  (.D(_02660_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .QN(_00644_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[528]$_DFFE_PN0P_  (.D(_02661_),
    .RN(net257),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .QN(_00675_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[529]$_DFFE_PN0P_  (.D(_02662_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .QN(_00706_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[52]$_DFFE_PN0P_  (.D(_02663_),
    .RN(net257),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .QN(_00784_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[530]$_DFFE_PN0P_  (.D(_02664_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .QN(_00737_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[531]$_DFFE_PN0P_  (.D(_02665_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .QN(_00768_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[532]$_DFFE_PN0P_  (.D(_02666_),
    .RN(net260),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .QN(_00799_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[533]$_DFFE_PN0P_  (.D(_02667_),
    .RN(net260),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .QN(_00830_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[534]$_DFFE_PN0P_  (.D(_02668_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .QN(_00861_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[535]$_DFFE_PN0P_  (.D(_02669_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .QN(_00892_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[536]$_DFFE_PN0P_  (.D(_02670_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .QN(_00923_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[537]$_DFFE_PN0P_  (.D(_02671_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .QN(_00954_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[538]$_DFFE_PN0P_  (.D(_02672_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .QN(_00985_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[539]$_DFFE_PN0P_  (.D(_02673_),
    .RN(net258),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .QN(_01016_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[53]$_DFFE_PN0P_  (.D(_02674_),
    .RN(net260),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .QN(_00815_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[540]$_DFFE_PN0P_  (.D(_02675_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .QN(_01047_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[541]$_DFFE_PN0P_  (.D(_02676_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .QN(_01078_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[542]$_DFFE_PN0P_  (.D(_02677_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .QN(_01109_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[543]$_DFFE_PN0P_  (.D(_02678_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .QN(_01140_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[544]$_DFFE_PN0P_  (.D(_02679_),
    .RN(net259),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .QN(_00202_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[545]$_DFFE_PN0P_  (.D(_02680_),
    .RN(net259),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .QN(_00157_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[546]$_DFFE_PN0P_  (.D(_02681_),
    .RN(net259),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .QN(_00264_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[547]$_DFFE_PN0P_  (.D(_02682_),
    .RN(net260),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .QN(_00295_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[548]$_DFFE_PN0P_  (.D(_02683_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .QN(_00325_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[549]$_DFFE_PN0P_  (.D(_02684_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .QN(_00355_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[54]$_DFFE_PN0P_  (.D(_02685_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .QN(_00846_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[550]$_DFFE_PN0P_  (.D(_02686_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .QN(_00385_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[551]$_DFFE_PN0P_  (.D(_02687_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .QN(_00415_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[552]$_DFFE_PN0P_  (.D(_02688_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .QN(_00445_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[553]$_DFFE_PN0P_  (.D(_02689_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .QN(_00475_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[554]$_DFFE_PN0P_  (.D(_02690_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .QN(_00505_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[555]$_DFFE_PN0P_  (.D(_02691_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .QN(_00535_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[556]$_DFFE_PN0P_  (.D(_02692_),
    .RN(net259),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .QN(_00234_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[557]$_DFFE_PN0P_  (.D(_02693_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .QN(_00583_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[558]$_DFFE_PN0P_  (.D(_02694_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .QN(_00614_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[559]$_DFFE_PN0P_  (.D(_02695_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .QN(_00645_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[55]$_DFFE_PN0P_  (.D(_02696_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .QN(_00877_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[560]$_DFFE_PN0P_  (.D(_02697_),
    .RN(net257),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .QN(_00676_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[561]$_DFFE_PN0P_  (.D(_02698_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .QN(_00707_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[562]$_DFFE_PN0P_  (.D(_02699_),
    .RN(net257),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .QN(_00738_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[563]$_DFFE_PN0P_  (.D(_02700_),
    .RN(net260),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .QN(_00769_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[564]$_DFFE_PN0P_  (.D(_02701_),
    .RN(net260),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .QN(_00800_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[565]$_DFFE_PN0P_  (.D(_02702_),
    .RN(net258),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .QN(_00831_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[566]$_DFFE_PN0P_  (.D(_02703_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .QN(_00862_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[567]$_DFFE_PN0P_  (.D(_02704_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .QN(_00893_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[568]$_DFFE_PN0P_  (.D(_02705_),
    .RN(net260),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .QN(_00924_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[569]$_DFFE_PN0P_  (.D(_02706_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .QN(_00955_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[56]$_DFFE_PN0P_  (.D(_02707_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .QN(_00908_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[570]$_DFFE_PN0P_  (.D(_02708_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .QN(_00986_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[571]$_DFFE_PN0P_  (.D(_02709_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .QN(_01017_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[572]$_DFFE_PN0P_  (.D(_02710_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .QN(_01048_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[573]$_DFFE_PN0P_  (.D(_02711_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .QN(_01079_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[574]$_DFFE_PN0P_  (.D(_02712_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .QN(_01110_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[575]$_DFFE_PN0P_  (.D(_02713_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .QN(_01141_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[576]$_DFFE_PN0P_  (.D(_02714_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .QN(_00203_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[577]$_DFFE_PN0P_  (.D(_02715_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .QN(_00158_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[578]$_DFFE_PN0P_  (.D(_02716_),
    .RN(net260),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .QN(_00265_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[579]$_DFFE_PN0P_  (.D(_02717_),
    .RN(net260),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .QN(_00296_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[57]$_DFFE_PN0P_  (.D(_02718_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .QN(_00939_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[580]$_DFFE_PN0P_  (.D(_02719_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .QN(_00326_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[581]$_DFFE_PN0P_  (.D(_02720_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .QN(_00356_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[582]$_DFFE_PN0P_  (.D(_02721_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .QN(_00386_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[583]$_DFFE_PN0P_  (.D(_02722_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .QN(_00416_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[584]$_DFFE_PN0P_  (.D(_02723_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .QN(_00446_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[585]$_DFFE_PN0P_  (.D(_02724_),
    .RN(net256),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .QN(_00476_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[586]$_DFFE_PN0P_  (.D(_02725_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .QN(_00506_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[587]$_DFFE_PN0P_  (.D(_02726_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .QN(_00536_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[588]$_DFFE_PN0P_  (.D(_02727_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .QN(_00235_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[589]$_DFFE_PN0P_  (.D(_02728_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .QN(_00584_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[58]$_DFFE_PN0P_  (.D(_02729_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .QN(_00970_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[590]$_DFFE_PN0P_  (.D(_02730_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .QN(_00615_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[591]$_DFFE_PN0P_  (.D(_02731_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .QN(_00646_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[592]$_DFFE_PN0P_  (.D(_02732_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .QN(_00677_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[593]$_DFFE_PN0P_  (.D(_02733_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .QN(_00708_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[594]$_DFFE_PN0P_  (.D(_02734_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .QN(_00739_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[595]$_DFFE_PN0P_  (.D(_02735_),
    .RN(net260),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .QN(_00770_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[596]$_DFFE_PN0P_  (.D(_02736_),
    .RN(net257),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .QN(_00801_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[597]$_DFFE_PN0P_  (.D(_02737_),
    .RN(net260),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .QN(_00832_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[598]$_DFFE_PN0P_  (.D(_02738_),
    .RN(net255),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .QN(_00863_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[599]$_DFFE_PN0P_  (.D(_02739_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .QN(_00894_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[59]$_DFFE_PN0P_  (.D(_02740_),
    .RN(net260),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .QN(_01001_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[5]$_DFFE_PN0P_  (.D(_02741_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .QN(_13620_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[600]$_DFFE_PN0P_  (.D(_02742_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .QN(_00925_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[601]$_DFFE_PN0P_  (.D(_02743_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .QN(_00956_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[602]$_DFFE_PN0P_  (.D(_02744_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .QN(_00987_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[603]$_DFFE_PN0P_  (.D(_02745_),
    .RN(net258),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .QN(_01018_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[604]$_DFFE_PN0P_  (.D(_02746_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .QN(_01049_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[605]$_DFFE_PN0P_  (.D(_02747_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .QN(_01080_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[606]$_DFFE_PN0P_  (.D(_02748_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .QN(_01111_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[607]$_DFFE_PN0P_  (.D(_02749_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .QN(_01142_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[608]$_DFFE_PN0P_  (.D(_02750_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .QN(_00204_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[609]$_DFFE_PN0P_  (.D(_02751_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .QN(_00159_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[60]$_DFFE_PN0P_  (.D(_02752_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .QN(_01032_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[610]$_DFFE_PN0P_  (.D(_02753_),
    .RN(net255),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .QN(_00266_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[611]$_DFFE_PN0P_  (.D(_02754_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .QN(_00297_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[612]$_DFFE_PN0P_  (.D(_02755_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .QN(_00327_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[613]$_DFFE_PN0P_  (.D(_02756_),
    .RN(net259),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .QN(_00357_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[614]$_DFFE_PN0P_  (.D(_02757_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .QN(_00387_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[615]$_DFFE_PN0P_  (.D(_02758_),
    .RN(net263),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .QN(_00417_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[616]$_DFFE_PN0P_  (.D(_02759_),
    .RN(net255),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .QN(_00447_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[617]$_DFFE_PN0P_  (.D(_02760_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .QN(_00477_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[618]$_DFFE_PN0P_  (.D(_02761_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .QN(_00507_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[619]$_DFFE_PN0P_  (.D(_02762_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .QN(_00537_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[61]$_DFFE_PN0P_  (.D(_02763_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .QN(_01063_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[620]$_DFFE_PN0P_  (.D(_02764_),
    .RN(net259),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .QN(_00236_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[621]$_DFFE_PN0P_  (.D(_02765_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .QN(_00585_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[622]$_DFFE_PN0P_  (.D(_02766_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .QN(_00616_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[623]$_DFFE_PN0P_  (.D(_02767_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .QN(_00647_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[624]$_DFFE_PN0P_  (.D(_02768_),
    .RN(net257),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .QN(_00678_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[625]$_DFFE_PN0P_  (.D(_02769_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .QN(_00709_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[626]$_DFFE_PN0P_  (.D(_02770_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .QN(_00740_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[627]$_DFFE_PN0P_  (.D(_02771_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .QN(_00771_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[628]$_DFFE_PN0P_  (.D(_02772_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .QN(_00802_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[629]$_DFFE_PN0P_  (.D(_02773_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .QN(_00833_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[62]$_DFFE_PN0P_  (.D(_02774_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .QN(_01094_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[630]$_DFFE_PN0P_  (.D(_02775_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .QN(_00864_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[631]$_DFFE_PN0P_  (.D(_02776_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .QN(_00895_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[632]$_DFFE_PN0P_  (.D(_02777_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .QN(_00926_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[633]$_DFFE_PN0P_  (.D(_02778_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .QN(_00957_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[634]$_DFFE_PN0P_  (.D(_02779_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .QN(_00988_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[635]$_DFFE_PN0P_  (.D(_02780_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .QN(_01019_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[636]$_DFFE_PN0P_  (.D(_02781_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .QN(_01050_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[637]$_DFFE_PN0P_  (.D(_02782_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .QN(_01081_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[638]$_DFFE_PN0P_  (.D(_02783_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .QN(_01112_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[639]$_DFFE_PN0P_  (.D(_02784_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .QN(_01143_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[63]$_DFFE_PN0P_  (.D(_02785_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .QN(_01125_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[640]$_DFFE_PN0P_  (.D(_02786_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .QN(_00205_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[641]$_DFFE_PN0P_  (.D(_02787_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .QN(_00160_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[642]$_DFFE_PN0P_  (.D(_02788_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .QN(_00267_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[643]$_DFFE_PN0P_  (.D(_02789_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .QN(_00298_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[644]$_DFFE_PN0P_  (.D(_02790_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .QN(_00328_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[645]$_DFFE_PN0P_  (.D(_02791_),
    .RN(net259),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .QN(_00358_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[646]$_DFFE_PN0P_  (.D(_02792_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .QN(_00388_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[647]$_DFFE_PN0P_  (.D(_02793_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .QN(_00418_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[648]$_DFFE_PN0P_  (.D(_02794_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .QN(_00448_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[649]$_DFFE_PN0P_  (.D(_02795_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .QN(_00478_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[64]$_DFFE_PN0P_  (.D(_02796_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .QN(_00187_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[650]$_DFFE_PN0P_  (.D(_02797_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .QN(_00508_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[651]$_DFFE_PN0P_  (.D(_02798_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .QN(_00538_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[652]$_DFFE_PN0P_  (.D(_02799_),
    .RN(net259),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .QN(_00237_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[653]$_DFFE_PN0P_  (.D(_02800_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .QN(_00586_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[654]$_DFFE_PN0P_  (.D(_02801_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .QN(_00617_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[655]$_DFFE_PN0P_  (.D(_02802_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .QN(_00648_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[656]$_DFFE_PN0P_  (.D(_02803_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .QN(_00679_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[657]$_DFFE_PN0P_  (.D(_02804_),
    .RN(net257),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .QN(_00710_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[658]$_DFFE_PN0P_  (.D(_02805_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .QN(_00741_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[659]$_DFFE_PN0P_  (.D(_02806_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .QN(_00772_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[65]$_DFFE_PN0P_  (.D(_02807_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .QN(_00142_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[660]$_DFFE_PN0P_  (.D(_02808_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .QN(_00803_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[661]$_DFFE_PN0P_  (.D(_02809_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .QN(_00834_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[662]$_DFFE_PN0P_  (.D(_02810_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .QN(_00865_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[663]$_DFFE_PN0P_  (.D(_02811_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .QN(_00896_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[664]$_DFFE_PN0P_  (.D(_02812_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .QN(_00927_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[665]$_DFFE_PN0P_  (.D(_02813_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .QN(_00958_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[666]$_DFFE_PN0P_  (.D(_02814_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .QN(_00989_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[667]$_DFFE_PN0P_  (.D(_02815_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .QN(_01020_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[668]$_DFFE_PN0P_  (.D(_02816_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .QN(_01051_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[669]$_DFFE_PN0P_  (.D(_02817_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .QN(_01082_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[66]$_DFFE_PN0P_  (.D(_02818_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .QN(_00249_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[670]$_DFFE_PN0P_  (.D(_02819_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .QN(_01113_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[671]$_DFFE_PN0P_  (.D(_02820_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .QN(_01144_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[672]$_DFFE_PN0P_  (.D(_02821_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .QN(_00206_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[673]$_DFFE_PN0P_  (.D(_02822_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .QN(_00161_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[674]$_DFFE_PN0P_  (.D(_02823_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .QN(_00268_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[675]$_DFFE_PN0P_  (.D(_02824_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .QN(_00299_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[676]$_DFFE_PN0P_  (.D(_02825_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .QN(_00329_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[677]$_DFFE_PN0P_  (.D(_02826_),
    .RN(net259),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .QN(_00359_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[678]$_DFFE_PN0P_  (.D(_02827_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .QN(_00389_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[679]$_DFFE_PN0P_  (.D(_02828_),
    .RN(net263),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .QN(_00419_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[67]$_DFFE_PN0P_  (.D(_02829_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .QN(_00280_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[680]$_DFFE_PN0P_  (.D(_02830_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .QN(_00449_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[681]$_DFFE_PN0P_  (.D(_02831_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .QN(_00479_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[682]$_DFFE_PN0P_  (.D(_02832_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .QN(_00509_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[683]$_DFFE_PN0P_  (.D(_02833_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .QN(_00539_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[684]$_DFFE_PN0P_  (.D(_02834_),
    .RN(net259),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .QN(_00238_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[685]$_DFFE_PN0P_  (.D(_02835_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .QN(_00587_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[686]$_DFFE_PN0P_  (.D(_02836_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .QN(_00618_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[687]$_DFFE_PN0P_  (.D(_02837_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .QN(_00649_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[688]$_DFFE_PN0P_  (.D(_02838_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .QN(_00680_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[689]$_DFFE_PN0P_  (.D(_02839_),
    .RN(net257),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .QN(_00711_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[68]$_DFFE_PN0P_  (.D(_02840_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .QN(_00310_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[690]$_DFFE_PN0P_  (.D(_02841_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .QN(_00742_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[691]$_DFFE_PN0P_  (.D(_02842_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .QN(_00773_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[692]$_DFFE_PN0P_  (.D(_02843_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .QN(_00804_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[693]$_DFFE_PN0P_  (.D(_02844_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .QN(_00835_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[694]$_DFFE_PN0P_  (.D(_02845_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .QN(_00866_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[695]$_DFFE_PN0P_  (.D(_02846_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .QN(_00897_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[696]$_DFFE_PN0P_  (.D(_02847_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .QN(_00928_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[697]$_DFFE_PN0P_  (.D(_02848_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .QN(_00959_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[698]$_DFFE_PN0P_  (.D(_02849_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .QN(_00990_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[699]$_DFFE_PN0P_  (.D(_02850_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .QN(_01021_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[69]$_DFFE_PN0P_  (.D(_02851_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .QN(_00340_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[6]$_DFFE_PN0P_  (.D(_02852_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .QN(_13619_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[700]$_DFFE_PN0P_  (.D(_02853_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .QN(_01052_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[701]$_DFFE_PN0P_  (.D(_02854_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .QN(_01083_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[702]$_DFFE_PN0P_  (.D(_02855_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .QN(_01114_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[703]$_DFFE_PN0P_  (.D(_02856_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .QN(_01145_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[704]$_DFFE_PN0P_  (.D(_02857_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .QN(_00207_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[705]$_DFFE_PN0P_  (.D(_02858_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .QN(_00162_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[706]$_DFFE_PN0P_  (.D(_02859_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .QN(_00269_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[707]$_DFFE_PN0P_  (.D(_02860_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .QN(_00300_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[708]$_DFFE_PN0P_  (.D(_02861_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .QN(_00330_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[709]$_DFFE_PN0P_  (.D(_02862_),
    .RN(net256),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .QN(_00360_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[70]$_DFFE_PN0P_  (.D(_02863_),
    .RN(net256),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .QN(_00370_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[710]$_DFFE_PN0P_  (.D(_02864_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .QN(_00390_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[711]$_DFFE_PN0P_  (.D(_02865_),
    .RN(net263),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .QN(_00420_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[712]$_DFFE_PN0P_  (.D(_02866_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .QN(_00450_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[713]$_DFFE_PN0P_  (.D(_02867_),
    .RN(net263),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .QN(_00480_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[714]$_DFFE_PN0P_  (.D(_02868_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .QN(_00510_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[715]$_DFFE_PN0P_  (.D(_02869_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .QN(_00540_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[716]$_DFFE_PN0P_  (.D(_02870_),
    .RN(net259),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .QN(_00239_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[717]$_DFFE_PN0P_  (.D(_02871_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .QN(_00588_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[718]$_DFFE_PN0P_  (.D(_02872_),
    .RN(net257),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .QN(_00619_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[719]$_DFFE_PN0P_  (.D(_02873_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .QN(_00650_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[71]$_DFFE_PN0P_  (.D(_02874_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .QN(_00400_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[720]$_DFFE_PN0P_  (.D(_02875_),
    .RN(net257),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .QN(_00681_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[721]$_DFFE_PN0P_  (.D(_02876_),
    .RN(net257),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .QN(_00712_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[722]$_DFFE_PN0P_  (.D(_02877_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .QN(_00743_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[723]$_DFFE_PN0P_  (.D(_02878_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .QN(_00774_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[724]$_DFFE_PN0P_  (.D(_02879_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .QN(_00805_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[725]$_DFFE_PN0P_  (.D(_02880_),
    .RN(net258),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .QN(_00836_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[726]$_DFFE_PN0P_  (.D(_02881_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .QN(_00867_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[727]$_DFFE_PN0P_  (.D(_02882_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .QN(_00898_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[728]$_DFFE_PN0P_  (.D(_02883_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .QN(_00929_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[729]$_DFFE_PN0P_  (.D(_02884_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .QN(_00960_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[72]$_DFFE_PN0P_  (.D(_02885_),
    .RN(net259),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .QN(_00430_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[730]$_DFFE_PN0P_  (.D(_02886_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .QN(_00991_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[731]$_DFFE_PN0P_  (.D(_02887_),
    .RN(net258),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .QN(_01022_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[732]$_DFFE_PN0P_  (.D(_02888_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .QN(_01053_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[733]$_DFFE_PN0P_  (.D(_02889_),
    .RN(net255),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .QN(_01084_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[734]$_DFFE_PN0P_  (.D(_02890_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .QN(_01115_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[735]$_DFFE_PN0P_  (.D(_02891_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .QN(_01146_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[736]$_DFFE_PN0P_  (.D(_02892_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .QN(_00208_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[737]$_DFFE_PN0P_  (.D(_02893_),
    .RN(net259),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .QN(_00163_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[738]$_DFFE_PN0P_  (.D(_02894_),
    .RN(net255),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .QN(_00270_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[739]$_DFFE_PN0P_  (.D(_02895_),
    .RN(net255),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .QN(_00301_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[73]$_DFFE_PN0P_  (.D(_02896_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .QN(_00460_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[740]$_DFFE_PN0P_  (.D(_02897_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .QN(_00331_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[741]$_DFFE_PN0P_  (.D(_02898_),
    .RN(net256),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .QN(_00361_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[742]$_DFFE_PN0P_  (.D(_02899_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .QN(_00391_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[743]$_DFFE_PN0P_  (.D(_02900_),
    .RN(net263),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .QN(_00421_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[744]$_DFFE_PN0P_  (.D(_02901_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .QN(_00451_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[745]$_DFFE_PN0P_  (.D(_02902_),
    .RN(net263),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .QN(_00481_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[746]$_DFFE_PN0P_  (.D(_02903_),
    .RN(net256),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .QN(_00511_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[747]$_DFFE_PN0P_  (.D(_02904_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .QN(_00541_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[748]$_DFFE_PN0P_  (.D(_02905_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .QN(_00240_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[749]$_DFFE_PN0P_  (.D(_02906_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .QN(_00589_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[74]$_DFFE_PN0P_  (.D(_02907_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .QN(_00490_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[750]$_DFFE_PN0P_  (.D(_02908_),
    .RN(net257),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .QN(_00620_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[751]$_DFFE_PN0P_  (.D(_02909_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .QN(_00651_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[752]$_DFFE_PN0P_  (.D(_02910_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .QN(_00682_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[753]$_DFFE_PN0P_  (.D(_02911_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .QN(_00713_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[754]$_DFFE_PN0P_  (.D(_02912_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .QN(_00744_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[755]$_DFFE_PN0P_  (.D(_02913_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .QN(_00775_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[756]$_DFFE_PN0P_  (.D(_02914_),
    .RN(net260),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .QN(_00806_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[757]$_DFFE_PN0P_  (.D(_02915_),
    .RN(net260),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .QN(_00837_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[758]$_DFFE_PN0P_  (.D(_02916_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .QN(_00868_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[759]$_DFFE_PN0P_  (.D(_02917_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .QN(_00899_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[75]$_DFFE_PN0P_  (.D(_02918_),
    .RN(net263),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .QN(_00520_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[760]$_DFFE_PN0P_  (.D(_02919_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .QN(_00930_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[761]$_DFFE_PN0P_  (.D(_02920_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .QN(_00961_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[762]$_DFFE_PN0P_  (.D(_02921_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .QN(_00992_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[763]$_DFFE_PN0P_  (.D(_02922_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .QN(_01023_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[764]$_DFFE_PN0P_  (.D(_02923_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .QN(_01054_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[765]$_DFFE_PN0P_  (.D(_02924_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .QN(_01085_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[766]$_DFFE_PN0P_  (.D(_02925_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .QN(_01116_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[767]$_DFFE_PN0P_  (.D(_02926_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .QN(_01147_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[768]$_DFFE_PN0P_  (.D(_02927_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .QN(_00209_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[769]$_DFFE_PN0P_  (.D(_02928_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .QN(_00164_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[76]$_DFFE_PN0P_  (.D(_02929_),
    .RN(net256),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .QN(_00219_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[770]$_DFFE_PN0P_  (.D(_02930_),
    .RN(net255),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .QN(_00271_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[771]$_DFFE_PN0P_  (.D(_02931_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .QN(_00302_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[772]$_DFFE_PN0P_  (.D(_02932_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .QN(_00332_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[773]$_DFFE_PN0P_  (.D(_02933_),
    .RN(net256),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .QN(_00362_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[774]$_DFFE_PN0P_  (.D(_02934_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .QN(_00392_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[775]$_DFFE_PN0P_  (.D(_02935_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .QN(_00422_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[776]$_DFFE_PN0P_  (.D(_02936_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .QN(_00452_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[777]$_DFFE_PN0P_  (.D(_02937_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .QN(_00482_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[778]$_DFFE_PN0P_  (.D(_02938_),
    .RN(net256),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .QN(_00512_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[779]$_DFFE_PN0P_  (.D(_02939_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .QN(_00542_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[77]$_DFFE_PN0P_  (.D(_02940_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .QN(_00568_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[780]$_DFFE_PN0P_  (.D(_02941_),
    .RN(net256),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .QN(_00241_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[781]$_DFFE_PN0P_  (.D(_02942_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .QN(_00590_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[782]$_DFFE_PN0P_  (.D(_02943_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .QN(_00621_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[783]$_DFFE_PN0P_  (.D(_02944_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .QN(_00652_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[784]$_DFFE_PN0P_  (.D(_02945_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .QN(_00683_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[785]$_DFFE_PN0P_  (.D(_02946_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .QN(_00714_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[786]$_DFFE_PN0P_  (.D(_02947_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .QN(_00745_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[787]$_DFFE_PN0P_  (.D(_02948_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .QN(_00776_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[788]$_DFFE_PN0P_  (.D(_02949_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .QN(_00807_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[789]$_DFFE_PN0P_  (.D(_02950_),
    .RN(net260),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .QN(_00838_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[78]$_DFFE_PN0P_  (.D(_02951_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .QN(_00599_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[790]$_DFFE_PN0P_  (.D(_02952_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .QN(_00869_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[791]$_DFFE_PN0P_  (.D(_02953_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .QN(_00900_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[792]$_DFFE_PN0P_  (.D(_02954_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .QN(_00931_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[793]$_DFFE_PN0P_  (.D(_02955_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .QN(_00962_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[794]$_DFFE_PN0P_  (.D(_02956_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .QN(_00993_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[795]$_DFFE_PN0P_  (.D(_02957_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .QN(_01024_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[796]$_DFFE_PN0P_  (.D(_02958_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .QN(_01055_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[797]$_DFFE_PN0P_  (.D(_02959_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .QN(_01086_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[798]$_DFFE_PN0P_  (.D(_02960_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .QN(_01117_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[799]$_DFFE_PN0P_  (.D(_02961_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .QN(_01148_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[79]$_DFFE_PN0P_  (.D(_02962_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .QN(_00630_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[7]$_DFFE_PN0P_  (.D(_02963_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .QN(_13618_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[800]$_DFFE_PN0P_  (.D(_02964_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .QN(_00210_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[801]$_DFFE_PN0P_  (.D(_02965_),
    .RN(net259),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .QN(_00165_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[802]$_DFFE_PN0P_  (.D(_02966_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .QN(_00272_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[803]$_DFFE_PN0P_  (.D(_02967_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .QN(_00303_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[804]$_DFFE_PN0P_  (.D(_02968_),
    .RN(net263),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .QN(_00333_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[805]$_DFFE_PN0P_  (.D(_02969_),
    .RN(net256),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .QN(_00363_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[806]$_DFFE_PN0P_  (.D(_02970_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .QN(_00393_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[807]$_DFFE_PN0P_  (.D(_02971_),
    .RN(net263),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .QN(_00423_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[808]$_DFFE_PN0P_  (.D(_02972_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .QN(_00453_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[809]$_DFFE_PN0P_  (.D(_02973_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .QN(_00483_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[80]$_DFFE_PN0P_  (.D(_02974_),
    .RN(net257),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .QN(_00661_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[810]$_DFFE_PN0P_  (.D(_02975_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .QN(_00513_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[811]$_DFFE_PN0P_  (.D(_02976_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .QN(_00543_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[812]$_DFFE_PN0P_  (.D(_02977_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .QN(_00242_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[813]$_DFFE_PN0P_  (.D(_02978_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .QN(_00591_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[814]$_DFFE_PN0P_  (.D(_02979_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .QN(_00622_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[815]$_DFFE_PN0P_  (.D(_02980_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .QN(_00653_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[816]$_DFFE_PN0P_  (.D(_02981_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .QN(_00684_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[817]$_DFFE_PN0P_  (.D(_02982_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .QN(_00715_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[818]$_DFFE_PN0P_  (.D(_02983_),
    .RN(net257),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .QN(_00746_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[819]$_DFFE_PN0P_  (.D(_02984_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .QN(_00777_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[81]$_DFFE_PN0P_  (.D(_02985_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .QN(_00692_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[820]$_DFFE_PN0P_  (.D(_02986_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .QN(_00808_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[821]$_DFFE_PN0P_  (.D(_02987_),
    .RN(net260),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .QN(_00839_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[822]$_DFFE_PN0P_  (.D(_02988_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .QN(_00870_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[823]$_DFFE_PN0P_  (.D(_02989_),
    .RN(net255),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .QN(_00901_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[824]$_DFFE_PN0P_  (.D(_02990_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .QN(_00932_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[825]$_DFFE_PN0P_  (.D(_02991_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .QN(_00963_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[826]$_DFFE_PN0P_  (.D(_02992_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .QN(_00994_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[827]$_DFFE_PN0P_  (.D(_02993_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .QN(_01025_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[828]$_DFFE_PN0P_  (.D(_02994_),
    .RN(net255),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .QN(_01056_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[829]$_DFFE_PN0P_  (.D(_02995_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .QN(_01087_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[82]$_DFFE_PN0P_  (.D(_02996_),
    .RN(net256),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .QN(_00723_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[830]$_DFFE_PN0P_  (.D(_02997_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .QN(_01118_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[831]$_DFFE_PN0P_  (.D(_02998_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .QN(_01149_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[832]$_DFFE_PN0P_  (.D(_02999_),
    .RN(net259),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .QN(_00211_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[833]$_DFFE_PN0P_  (.D(_03000_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .QN(_00166_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[834]$_DFFE_PN0P_  (.D(_03001_),
    .RN(net255),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .QN(_00273_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[835]$_DFFE_PN0P_  (.D(_03002_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .QN(_00304_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[836]$_DFFE_PN0P_  (.D(_03003_),
    .RN(net263),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .QN(_00334_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[837]$_DFFE_PN0P_  (.D(_03004_),
    .RN(net256),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .QN(_00364_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[838]$_DFFE_PN0P_  (.D(_03005_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .QN(_00394_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[839]$_DFFE_PN0P_  (.D(_03006_),
    .RN(net263),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .QN(_00424_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[83]$_DFFE_PN0P_  (.D(_03007_),
    .RN(net260),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .QN(_00754_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[840]$_DFFE_PN0P_  (.D(_03008_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .QN(_00454_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[841]$_DFFE_PN0P_  (.D(_03009_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .QN(_00484_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[842]$_DFFE_PN0P_  (.D(_03010_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .QN(_00514_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[843]$_DFFE_PN0P_  (.D(_03011_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .QN(_00544_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[844]$_DFFE_PN0P_  (.D(_03012_),
    .RN(net256),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .QN(_00243_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[845]$_DFFE_PN0P_  (.D(_03013_),
    .RN(net256),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .QN(_00592_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[846]$_DFFE_PN0P_  (.D(_03014_),
    .RN(net257),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .QN(_00623_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[847]$_DFFE_PN0P_  (.D(_03015_),
    .RN(net257),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .QN(_00654_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[848]$_DFFE_PN0P_  (.D(_03016_),
    .RN(net257),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .QN(_00685_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[849]$_DFFE_PN0P_  (.D(_03017_),
    .RN(net257),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .QN(_00716_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[84]$_DFFE_PN0P_  (.D(_03018_),
    .RN(net257),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .QN(_00785_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[850]$_DFFE_PN0P_  (.D(_03019_),
    .RN(net256),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .QN(_00747_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[851]$_DFFE_PN0P_  (.D(_03020_),
    .RN(net255),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .QN(_00778_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[852]$_DFFE_PN0P_  (.D(_03021_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .QN(_00809_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[853]$_DFFE_PN0P_  (.D(_03022_),
    .RN(net260),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .QN(_00840_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[854]$_DFFE_PN0P_  (.D(_03023_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .QN(_00871_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[855]$_DFFE_PN0P_  (.D(_03024_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .QN(_00902_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[856]$_DFFE_PN0P_  (.D(_03025_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .QN(_00933_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[857]$_DFFE_PN0P_  (.D(_03026_),
    .RN(net255),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .QN(_00964_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[858]$_DFFE_PN0P_  (.D(_03027_),
    .RN(net255),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .QN(_00995_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[859]$_DFFE_PN0P_  (.D(_03028_),
    .RN(net258),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .QN(_01026_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[85]$_DFFE_PN0P_  (.D(_03029_),
    .RN(net260),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .QN(_00816_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[860]$_DFFE_PN0P_  (.D(_03030_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .QN(_01057_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[861]$_DFFE_PN0P_  (.D(_03031_),
    .RN(net255),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .QN(_01088_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[862]$_DFFE_PN0P_  (.D(_03032_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .QN(_01119_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[863]$_DFFE_PN0P_  (.D(_03033_),
    .RN(net255),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .QN(_01150_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[864]$_DFFE_PN0P_  (.D(_03034_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .QN(_00212_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[865]$_DFFE_PN0P_  (.D(_03035_),
    .RN(net259),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .QN(_00167_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[866]$_DFFE_PN0P_  (.D(_03036_),
    .RN(net260),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .QN(_00274_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[867]$_DFFE_PN0P_  (.D(_03037_),
    .RN(net259),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .QN(_00305_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[868]$_DFFE_PN0P_  (.D(_03038_),
    .RN(net263),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .QN(_00335_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[869]$_DFFE_PN0P_  (.D(_03039_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .QN(_00365_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[86]$_DFFE_PN0P_  (.D(_03040_),
    .RN(net258),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .QN(_00847_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[870]$_DFFE_PN0P_  (.D(_03041_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .QN(_00395_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[871]$_DFFE_PN0P_  (.D(_03042_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .QN(_00425_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[872]$_DFFE_PN0P_  (.D(_03043_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .QN(_00455_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[873]$_DFFE_PN0P_  (.D(_03044_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .QN(_00485_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[874]$_DFFE_PN0P_  (.D(_03045_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .QN(_00515_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[875]$_DFFE_PN0P_  (.D(_03046_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .QN(_00545_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[876]$_DFFE_PN0P_  (.D(_03047_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .QN(_00244_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[877]$_DFFE_PN0P_  (.D(_03048_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .QN(_00593_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[878]$_DFFE_PN0P_  (.D(_03049_),
    .RN(net257),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .QN(_00624_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[879]$_DFFE_PN0P_  (.D(_03050_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .QN(_00655_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[87]$_DFFE_PN0P_  (.D(_03051_),
    .RN(net258),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .QN(_00878_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[880]$_DFFE_PN0P_  (.D(_03052_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .QN(_00686_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[881]$_DFFE_PN0P_  (.D(_03053_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .QN(_00717_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[882]$_DFFE_PN0P_  (.D(_03054_),
    .RN(net257),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .QN(_00748_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[883]$_DFFE_PN0P_  (.D(_03055_),
    .RN(net260),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .QN(_00779_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[884]$_DFFE_PN0P_  (.D(_03056_),
    .RN(net260),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .QN(_00810_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[885]$_DFFE_PN0P_  (.D(_03057_),
    .RN(net258),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .QN(_00841_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[886]$_DFFE_PN0P_  (.D(_03058_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .QN(_00872_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[887]$_DFFE_PN0P_  (.D(_03059_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .QN(_00903_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[888]$_DFFE_PN0P_  (.D(_03060_),
    .RN(net260),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .QN(_00934_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[889]$_DFFE_PN0P_  (.D(_03061_),
    .RN(net260),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .QN(_00965_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[88]$_DFFE_PN0P_  (.D(_03062_),
    .RN(net260),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .QN(_00909_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[890]$_DFFE_PN0P_  (.D(_03063_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .QN(_00996_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[891]$_DFFE_PN0P_  (.D(_03064_),
    .RN(net258),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .QN(_01027_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[892]$_DFFE_PN0P_  (.D(_03065_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .QN(_01058_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[893]$_DFFE_PN0P_  (.D(_03066_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .QN(_01089_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[894]$_DFFE_PN0P_  (.D(_03067_),
    .RN(net258),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .QN(_01120_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[895]$_DFFE_PN0P_  (.D(_03068_),
    .RN(net260),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .QN(_01151_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[896]$_DFFE_PN0P_  (.D(_03069_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .QN(_00213_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[897]$_DFFE_PN0P_  (.D(_03070_),
    .RN(net259),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .QN(_00168_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[898]$_DFFE_PN0P_  (.D(_03071_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .QN(_00275_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[899]$_DFFE_PN0P_  (.D(_03072_),
    .RN(net259),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .QN(_00306_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[89]$_DFFE_PN0P_  (.D(_03073_),
    .RN(net259),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .QN(_00940_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[8]$_DFFE_PN0P_  (.D(_03074_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .QN(_13617_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[900]$_DFFE_PN0P_  (.D(_03075_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .QN(_00336_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[901]$_DFFE_PN0P_  (.D(_03076_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .QN(_00366_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[902]$_DFFE_PN0P_  (.D(_03077_),
    .RN(net256),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .QN(_00396_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[903]$_DFFE_PN0P_  (.D(_03078_),
    .RN(net263),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .QN(_00426_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[904]$_DFFE_PN0P_  (.D(_03079_),
    .RN(net259),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .QN(_00456_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[905]$_DFFE_PN0P_  (.D(_03080_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .QN(_00486_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[906]$_DFFE_PN0P_  (.D(_03081_),
    .RN(net256),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .QN(_00516_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[907]$_DFFE_PN0P_  (.D(_03082_),
    .RN(net263),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .QN(_00546_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[908]$_DFFE_PN0P_  (.D(_03083_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .QN(_00245_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[909]$_DFFE_PN0P_  (.D(_03084_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .QN(_00594_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[90]$_DFFE_PN0P_  (.D(_03085_),
    .RN(net258),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .QN(_00971_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[910]$_DFFE_PN0P_  (.D(_03086_),
    .RN(net257),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .QN(_00625_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[911]$_DFFE_PN0P_  (.D(_03087_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .QN(_00656_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[912]$_DFFE_PN0P_  (.D(_03088_),
    .RN(net257),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .QN(_00687_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[913]$_DFFE_PN0P_  (.D(_03089_),
    .RN(net257),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .QN(_00718_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[914]$_DFFE_PN0P_  (.D(_03090_),
    .RN(net257),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .QN(_00749_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[915]$_DFFE_PN0P_  (.D(_03091_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .QN(_00780_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[916]$_DFFE_PN0P_  (.D(_03092_),
    .RN(net260),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .QN(_00811_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[917]$_DFFE_PN0P_  (.D(_01184_),
    .RN(net260),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .QN(_00842_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[918]$_DFFE_PN0P_  (.D(_01185_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .QN(_00873_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[919]$_DFFE_PN0P_  (.D(_01186_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .QN(_00904_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[91]$_DFFE_PN0P_  (.D(_01187_),
    .RN(net258),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .QN(_01002_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[920]$_DFFE_PN0P_  (.D(_01188_),
    .RN(net255),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .QN(_00935_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[921]$_DFFE_PN0P_  (.D(_01189_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .QN(_00966_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[922]$_DFFE_PN0P_  (.D(_01190_),
    .RN(net255),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .QN(_00997_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[923]$_DFFE_PN0P_  (.D(_01191_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .QN(_01028_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[924]$_DFFE_PN0P_  (.D(_01192_),
    .RN(net255),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .QN(_01059_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[925]$_DFFE_PN0P_  (.D(_01193_),
    .RN(net260),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .QN(_01090_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[926]$_DFFE_PN0P_  (.D(_01194_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .QN(_01121_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[927]$_DFFE_PN0P_  (.D(_01195_),
    .RN(net260),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .QN(_01152_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[928]$_DFFE_PN0P_  (.D(_01196_),
    .RN(net259),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .QN(_00214_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[929]$_DFFE_PN0P_  (.D(_01197_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .QN(_00169_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[92]$_DFFE_PN0P_  (.D(_01198_),
    .RN(net258),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .QN(_01033_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[930]$_DFFE_PN0P_  (.D(_01199_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .QN(_00276_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[931]$_DFFE_PN0P_  (.D(_01200_),
    .RN(net259),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .QN(_00307_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[932]$_DFFE_PN0P_  (.D(_01201_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .QN(_00337_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[933]$_DFFE_PN0P_  (.D(_01202_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .QN(_00367_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[934]$_DFFE_PN0P_  (.D(_01203_),
    .RN(net263),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .QN(_00397_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[935]$_DFFE_PN0P_  (.D(_01204_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .QN(_00427_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[936]$_DFFE_PN0P_  (.D(_01205_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .QN(_00457_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[937]$_DFFE_PN0P_  (.D(_01206_),
    .RN(net263),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .QN(_00487_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[938]$_DFFE_PN0P_  (.D(_01207_),
    .RN(net256),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .QN(_00517_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[939]$_DFFE_PN0P_  (.D(_01208_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .QN(_00547_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[93]$_DFFE_PN0P_  (.D(_01209_),
    .RN(net260),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .QN(_01064_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[940]$_DFFE_PN0P_  (.D(_01210_),
    .RN(net259),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .QN(_00246_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[941]$_DFFE_PN0P_  (.D(_01211_),
    .RN(net256),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .QN(_00595_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[942]$_DFFE_PN0P_  (.D(_01212_),
    .RN(net257),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .QN(_00626_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[943]$_DFFE_PN0P_  (.D(_01213_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .QN(_00657_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[944]$_DFFE_PN0P_  (.D(_01214_),
    .RN(net260),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .QN(_00688_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[945]$_DFFE_PN0P_  (.D(_01215_),
    .RN(net260),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .QN(_00719_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[946]$_DFFE_PN0P_  (.D(_01216_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .QN(_00750_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[947]$_DFFE_PN0P_  (.D(_01217_),
    .RN(net255),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .QN(_00781_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[948]$_DFFE_PN0P_  (.D(_01218_),
    .RN(net260),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .QN(_00812_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[949]$_DFFE_PN0P_  (.D(_01219_),
    .RN(net258),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .QN(_00843_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[94]$_DFFE_PN0P_  (.D(_01220_),
    .RN(net260),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .QN(_01095_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[950]$_DFFE_PN0P_  (.D(_01221_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .QN(_00874_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[951]$_DFFE_PN0P_  (.D(_01222_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .QN(_00905_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[952]$_DFFE_PN0P_  (.D(_01223_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .QN(_00936_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[953]$_DFFE_PN0P_  (.D(_01224_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .QN(_00967_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[954]$_DFFE_PN0P_  (.D(_01225_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .QN(_00998_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[955]$_DFFE_PN0P_  (.D(_01226_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .QN(_01029_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[956]$_DFFE_PN0P_  (.D(_01227_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .QN(_01060_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[957]$_DFFE_PN0P_  (.D(_01228_),
    .RN(net260),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .QN(_01091_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[958]$_DFFE_PN0P_  (.D(_01229_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .QN(_01122_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[959]$_DFFE_PN0P_  (.D(_01230_),
    .RN(net259),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .QN(_01153_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[95]$_DFFE_PN0P_  (.D(_01231_),
    .RN(net259),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .QN(_01126_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[960]$_DFFE_PN0P_  (.D(_01232_),
    .RN(net259),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .QN(_00215_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[961]$_DFFE_PN0P_  (.D(_01233_),
    .RN(net259),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .QN(_00170_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[962]$_DFFE_PN0P_  (.D(_01234_),
    .RN(net260),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .QN(_00277_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[963]$_DFFE_PN0P_  (.D(_01235_),
    .RN(net259),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .QN(_00308_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[964]$_DFFE_PN0P_  (.D(_01236_),
    .RN(net263),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .QN(_00338_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[965]$_DFFE_PN0P_  (.D(_01237_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .QN(_00368_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[966]$_DFFE_PN0P_  (.D(_01238_),
    .RN(net259),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .QN(_00398_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[967]$_DFFE_PN0P_  (.D(_01239_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .QN(_00428_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[968]$_DFFE_PN0P_  (.D(_01240_),
    .RN(net259),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .QN(_00458_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[969]$_DFFE_PN0P_  (.D(_01241_),
    .RN(net263),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .QN(_00488_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[96]$_DFFE_PN0P_  (.D(_01242_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .QN(_00188_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[970]$_DFFE_PN0P_  (.D(_01243_),
    .RN(net256),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .QN(_00518_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[971]$_DFFE_PN0P_  (.D(_01244_),
    .RN(net263),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .QN(_00548_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[972]$_DFFE_PN0P_  (.D(_01245_),
    .RN(net259),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .QN(_00247_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[973]$_DFFE_PN0P_  (.D(_01246_),
    .RN(net256),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .QN(_00596_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[974]$_DFFE_PN0P_  (.D(_01247_),
    .RN(net257),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .QN(_00627_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[975]$_DFFE_PN0P_  (.D(_01248_),
    .RN(net257),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .QN(_00658_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[976]$_DFFE_PN0P_  (.D(_01249_),
    .RN(net257),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .QN(_00689_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[977]$_DFFE_PN0P_  (.D(_01250_),
    .RN(net260),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .QN(_00720_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[978]$_DFFE_PN0P_  (.D(_01251_),
    .RN(net257),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .QN(_00751_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[979]$_DFFE_PN0P_  (.D(_01252_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .QN(_00782_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[97]$_DFFE_PN0P_  (.D(_01253_),
    .RN(net259),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .QN(_00143_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[980]$_DFFE_PN0P_  (.D(_01254_),
    .RN(net260),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .QN(_00813_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[981]$_DFFE_PN0P_  (.D(_01255_),
    .RN(net258),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .QN(_00844_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[982]$_DFFE_PN0P_  (.D(_01256_),
    .RN(net255),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .QN(_00875_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[983]$_DFFE_PN0P_  (.D(_01257_),
    .RN(net255),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .QN(_00906_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[984]$_DFFE_PN0P_  (.D(_01258_),
    .RN(net255),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .QN(_00937_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[985]$_DFFE_PN0P_  (.D(_01259_),
    .RN(net255),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .QN(_00968_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[986]$_DFFE_PN0P_  (.D(_01260_),
    .RN(net255),
    .CK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .QN(_00999_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[987]$_DFFE_PN0P_  (.D(_01261_),
    .RN(net258),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .QN(_01030_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[988]$_DFFE_PN0P_  (.D(_01262_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .QN(_01061_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[989]$_DFFE_PN0P_  (.D(_01263_),
    .RN(net260),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .QN(_01092_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[98]$_DFFE_PN0P_  (.D(_01264_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .QN(_00250_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[990]$_DFFE_PN0P_  (.D(_01265_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .QN(_01123_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[991]$_DFFE_PN0P_  (.D(_01266_),
    .RN(net260),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .QN(_01154_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[99]$_DFFE_PN0P_  (.D(_01267_),
    .RN(net259),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .QN(_00281_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[9]$_DFFE_PN0P_  (.D(_01268_),
    .RN(net256),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .QN(_13616_));
 DFFR_X2 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_01269_),
    .RN(net261),
    .CK(clknet_leaf_111_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .QN(_13615_));
 DFFR_X1 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_01270_),
    .RN(net261),
    .CK(clknet_leaf_111_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .QN(_13614_));
 DFFR_X1 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_01271_),
    .RN(net261),
    .CK(clknet_leaf_110_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .QN(_13613_));
 DFFR_X2 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_01272_),
    .RN(net261),
    .CK(clknet_leaf_110_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .QN(_13612_));
 DFFR_X1 \id_stage_i.controller_i.debug_mode_q$_DFFE_PN0P_  (.D(_01273_),
    .RN(net262),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.debug_mode_i ),
    .QN(_01156_));
 DFFR_X1 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .RN(net262),
    .CK(clknet_leaf_109_clk),
    .Q(\id_stage_i.controller_i.exc_req_q ),
    .QN(_14054_));
 DFFR_X1 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .RN(net262),
    .CK(clknet_leaf_109_clk),
    .Q(\id_stage_i.controller_i.illegal_insn_q ),
    .QN(_01157_));
 DFFR_X1 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_d ),
    .RN(net262),
    .CK(clknet_leaf_110_clk),
    .Q(\id_stage_i.controller_i.load_err_q ),
    .QN(_13611_));
 DFFR_X1 \id_stage_i.controller_i.nmi_mode_q$_DFFE_PN0P_  (.D(_01274_),
    .RN(net265),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.nmi_mode_i ),
    .QN(_14055_));
 DFFR_X1 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_d ),
    .RN(net262),
    .CK(clknet_leaf_109_clk),
    .Q(\id_stage_i.controller_i.store_err_q ),
    .QN(_14056_));
 DFFR_X1 \id_stage_i.g_branch_set_flop.branch_set_q$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .RN(net262),
    .CK(clknet_leaf_109_clk),
    .Q(\id_stage_i.branch_set ),
    .QN(_13610_));
 DFFR_X1 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_01275_),
    .RN(net261),
    .CK(clknet_leaf_111_clk),
    .Q(\id_stage_i.id_fsm_q ),
    .QN(_13609_));
 DFFR_X1 \id_stage_i.imd_val_q[0]$_DFFE_PN0P_  (.D(_01276_),
    .RN(net263),
    .CK(clknet_leaf_18_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .QN(_13608_));
 DFFR_X1 \id_stage_i.imd_val_q[10]$_DFFE_PN0P_  (.D(_01277_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .QN(_13607_));
 DFFR_X1 \id_stage_i.imd_val_q[11]$_DFFE_PN0P_  (.D(_01278_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .QN(_13606_));
 DFFR_X1 \id_stage_i.imd_val_q[12]$_DFFE_PN0P_  (.D(_01279_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .QN(_13605_));
 DFFR_X1 \id_stage_i.imd_val_q[13]$_DFFE_PN0P_  (.D(_01280_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .QN(_13604_));
 DFFR_X1 \id_stage_i.imd_val_q[14]$_DFFE_PN0P_  (.D(_01281_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .QN(_13603_));
 DFFR_X1 \id_stage_i.imd_val_q[15]$_DFFE_PN0P_  (.D(_01282_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .QN(_13602_));
 DFFR_X1 \id_stage_i.imd_val_q[16]$_DFFE_PN0P_  (.D(_01283_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .QN(_13601_));
 DFFR_X1 \id_stage_i.imd_val_q[17]$_DFFE_PN0P_  (.D(_01284_),
    .RN(net264),
    .CK(clknet_leaf_18_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .QN(_13600_));
 DFFR_X1 \id_stage_i.imd_val_q[18]$_DFFE_PN0P_  (.D(_01285_),
    .RN(net264),
    .CK(clknet_leaf_18_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .QN(_13599_));
 DFFR_X1 \id_stage_i.imd_val_q[19]$_DFFE_PN0P_  (.D(_01286_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .QN(_13598_));
 DFFR_X1 \id_stage_i.imd_val_q[1]$_DFFE_PN0P_  (.D(_01287_),
    .RN(net264),
    .CK(clknet_leaf_18_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .QN(_13597_));
 DFFR_X1 \id_stage_i.imd_val_q[20]$_DFFE_PN0P_  (.D(_01288_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .QN(_13596_));
 DFFR_X1 \id_stage_i.imd_val_q[21]$_DFFE_PN0P_  (.D(_01289_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .QN(_13595_));
 DFFR_X1 \id_stage_i.imd_val_q[22]$_DFFE_PN0P_  (.D(_01290_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .QN(_13594_));
 DFFR_X1 \id_stage_i.imd_val_q[23]$_DFFE_PN0P_  (.D(_01291_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .QN(_13593_));
 DFFR_X1 \id_stage_i.imd_val_q[24]$_DFFE_PN0P_  (.D(_01292_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .QN(_13592_));
 DFFR_X1 \id_stage_i.imd_val_q[25]$_DFFE_PN0P_  (.D(_01293_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .QN(_13591_));
 DFFR_X1 \id_stage_i.imd_val_q[26]$_DFFE_PN0P_  (.D(_01294_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .QN(_13590_));
 DFFR_X1 \id_stage_i.imd_val_q[27]$_DFFE_PN0P_  (.D(_01295_),
    .RN(net263),
    .CK(clknet_leaf_14_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .QN(_13589_));
 DFFR_X1 \id_stage_i.imd_val_q[28]$_DFFE_PN0P_  (.D(_01296_),
    .RN(net263),
    .CK(clknet_leaf_16_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .QN(_13588_));
 DFFR_X1 \id_stage_i.imd_val_q[29]$_DFFE_PN0P_  (.D(_01297_),
    .RN(net263),
    .CK(clknet_leaf_15_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .QN(_13587_));
 DFFR_X1 \id_stage_i.imd_val_q[2]$_DFFE_PN0P_  (.D(_01298_),
    .RN(net263),
    .CK(clknet_leaf_17_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .QN(_13586_));
 DFFR_X1 \id_stage_i.imd_val_q[30]$_DFFE_PN0P_  (.D(_01299_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .QN(_13585_));
 DFFR_X2 \id_stage_i.imd_val_q[31]$_DFFE_PN0P_  (.D(_01300_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .QN(_13584_));
 DFFR_X1 \id_stage_i.imd_val_q[34]$_DFFE_PN0P_  (.D(_01301_),
    .RN(net264),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .QN(_00217_));
 DFFR_X2 \id_stage_i.imd_val_q[35]$_DFFE_PN0P_  (.D(_01302_),
    .RN(net264),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .QN(_00185_));
 DFFR_X2 \id_stage_i.imd_val_q[36]$_DFFE_PN0P_  (.D(_01303_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .QN(_00556_));
 DFFR_X2 \id_stage_i.imd_val_q[37]$_DFFE_PN0P_  (.D(_01304_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .QN(_00557_));
 DFFR_X2 \id_stage_i.imd_val_q[38]$_DFFE_PN0P_  (.D(_01305_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .QN(_00558_));
 DFFR_X2 \id_stage_i.imd_val_q[39]$_DFFE_PN0P_  (.D(_01306_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .QN(_00559_));
 DFFR_X1 \id_stage_i.imd_val_q[3]$_DFFE_PN0P_  (.D(_01307_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .QN(_13583_));
 DFFR_X2 \id_stage_i.imd_val_q[40]$_DFFE_PN0P_  (.D(_01308_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .QN(_00560_));
 DFFR_X2 \id_stage_i.imd_val_q[41]$_DFFE_PN0P_  (.D(_01309_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .QN(_00561_));
 DFFR_X2 \id_stage_i.imd_val_q[42]$_DFFE_PN0P_  (.D(_01310_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .QN(_00562_));
 DFFR_X2 \id_stage_i.imd_val_q[43]$_DFFE_PN0P_  (.D(_01311_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .QN(_00563_));
 DFFR_X2 \id_stage_i.imd_val_q[44]$_DFFE_PN0P_  (.D(_01312_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .QN(_00564_));
 DFFR_X2 \id_stage_i.imd_val_q[45]$_DFFE_PN0P_  (.D(_01313_),
    .RN(net264),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .QN(_00565_));
 DFFR_X2 \id_stage_i.imd_val_q[46]$_DFFE_PN0P_  (.D(_01314_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .QN(_00566_));
 DFFR_X1 \id_stage_i.imd_val_q[47]$_DFFE_PN0P_  (.D(_01315_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .QN(_00597_));
 DFFR_X1 \id_stage_i.imd_val_q[48]$_DFFE_PN0P_  (.D(_01316_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .QN(_00628_));
 DFFR_X2 \id_stage_i.imd_val_q[49]$_DFFE_PN0P_  (.D(_01317_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .QN(_00659_));
 DFFR_X1 \id_stage_i.imd_val_q[4]$_DFFE_PN0P_  (.D(_01318_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .QN(_13582_));
 DFFR_X1 \id_stage_i.imd_val_q[50]$_DFFE_PN0P_  (.D(_01319_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .QN(_00690_));
 DFFR_X2 \id_stage_i.imd_val_q[51]$_DFFE_PN0P_  (.D(_01320_),
    .RN(net264),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .QN(_00721_));
 DFFR_X2 \id_stage_i.imd_val_q[52]$_DFFE_PN0P_  (.D(_01321_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .QN(_00752_));
 DFFR_X2 \id_stage_i.imd_val_q[53]$_DFFE_PN0P_  (.D(_01322_),
    .RN(net264),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .QN(_00783_));
 DFFR_X2 \id_stage_i.imd_val_q[54]$_DFFE_PN0P_  (.D(_01323_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .QN(_00814_));
 DFFR_X2 \id_stage_i.imd_val_q[55]$_DFFE_PN0P_  (.D(_01324_),
    .RN(net264),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .QN(_00845_));
 DFFR_X2 \id_stage_i.imd_val_q[56]$_DFFE_PN0P_  (.D(_01325_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .QN(_00876_));
 DFFR_X2 \id_stage_i.imd_val_q[57]$_DFFE_PN0P_  (.D(_01326_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .QN(_00907_));
 DFFR_X2 \id_stage_i.imd_val_q[58]$_DFFE_PN0P_  (.D(_01327_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .QN(_00938_));
 DFFR_X2 \id_stage_i.imd_val_q[59]$_DFFE_PN0P_  (.D(_01328_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .QN(_00969_));
 DFFR_X1 \id_stage_i.imd_val_q[5]$_DFFE_PN0P_  (.D(_01329_),
    .RN(net263),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .QN(_13581_));
 DFFR_X2 \id_stage_i.imd_val_q[60]$_DFFE_PN0P_  (.D(_01330_),
    .RN(net264),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .QN(_01000_));
 DFFR_X2 \id_stage_i.imd_val_q[61]$_DFFE_PN0P_  (.D(_01331_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .QN(_01031_));
 DFFR_X2 \id_stage_i.imd_val_q[62]$_DFFE_PN0P_  (.D(_01332_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .QN(_01062_));
 DFFR_X2 \id_stage_i.imd_val_q[63]$_DFFE_PN0P_  (.D(_01333_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .QN(_01093_));
 DFFR_X2 \id_stage_i.imd_val_q[64]$_DFFE_PN0P_  (.D(_01334_),
    .RN(net264),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .QN(_01124_));
 DFFR_X1 \id_stage_i.imd_val_q[65]$_DFFE_PN0P_  (.D(_01335_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .QN(_01155_));
 DFFR_X1 \id_stage_i.imd_val_q[66]$_DFFE_PN0P_  (.D(_01336_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .QN(_13580_));
 DFFR_X1 \id_stage_i.imd_val_q[67]$_DFFE_PN0P_  (.D(_01337_),
    .RN(net264),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .QN(_00132_));
 DFFR_X1 \id_stage_i.imd_val_q[6]$_DFFE_PN0P_  (.D(_01338_),
    .RN(net263),
    .CK(clknet_leaf_20_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .QN(_13579_));
 DFFR_X1 \id_stage_i.imd_val_q[7]$_DFFE_PN0P_  (.D(_01339_),
    .RN(net263),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .QN(_13578_));
 DFFR_X1 \id_stage_i.imd_val_q[8]$_DFFE_PN0P_  (.D(_01340_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .QN(_13577_));
 DFFR_X1 \id_stage_i.imd_val_q[9]$_DFFE_PN0P_  (.D(_01341_),
    .RN(net263),
    .CK(clknet_leaf_19_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .QN(_14057_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .RN(net261),
    .CK(clknet_leaf_114_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .QN(_14058_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .RN(net261),
    .CK(clknet_leaf_114_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .QN(_14059_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .RN(net261),
    .CK(clknet_leaf_110_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .QN(_13576_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(_01342_),
    .CK(clknet_leaf_39_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .QN(_13575_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(_01343_),
    .CK(clknet_leaf_43_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .QN(_13574_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(_01344_),
    .CK(clknet_leaf_43_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .QN(_13573_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(_01345_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .QN(_13572_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(_01346_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .QN(_13571_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(_01347_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .QN(_13570_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(_01348_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .QN(_13569_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(_01349_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .QN(_13568_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(_01350_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .QN(_13567_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(_01351_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .QN(_13566_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(_01352_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .QN(_13565_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(_01353_),
    .CK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .QN(_13564_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(_01354_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .QN(_13563_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(_01355_),
    .CK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .QN(_13562_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(_01356_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .QN(_13561_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(_01357_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .QN(_13560_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(_01358_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .QN(_13559_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(_01359_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .QN(_13558_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(_01360_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .QN(_13557_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(_01361_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .QN(_13556_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(_01362_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .QN(_13555_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(_01363_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .QN(_13554_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(_01364_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .QN(_13553_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(_01365_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .QN(_13552_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(_01366_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .QN(_13551_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(_01367_),
    .CK(clknet_leaf_43_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .QN(_13550_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(_01368_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .QN(_13549_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(_01369_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .QN(_13548_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(_01370_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .QN(_13547_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(_01371_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .QN(_13546_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(_01372_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .QN(_13545_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(_01373_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .QN(_13544_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(_01374_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .QN(_13543_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(_01375_),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.pc_if_i[1] ),
    .QN(_00137_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(_01376_),
    .CK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.pc_if_i[11] ),
    .QN(_13542_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(_01377_),
    .CK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.pc_if_i[12] ),
    .QN(_13541_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(_01378_),
    .CK(clknet_leaf_43_clk),
    .Q(\cs_registers_i.pc_if_i[13] ),
    .QN(_13540_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(_01379_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[14] ),
    .QN(_13539_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(_01380_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[15] ),
    .QN(_13538_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(_01381_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[16] ),
    .QN(_13537_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(_01382_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_if_i[17] ),
    .QN(_13536_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(_01383_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[18] ),
    .QN(_13535_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(_01384_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_if_i[19] ),
    .QN(_13534_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(_01385_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[20] ),
    .QN(_13533_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(_01386_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[2] ),
    .QN(_15352_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(_01387_),
    .CK(clknet_leaf_39_clk),
    .Q(\cs_registers_i.pc_if_i[21] ),
    .QN(_13532_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(_01388_),
    .CK(clknet_leaf_43_clk),
    .Q(\cs_registers_i.pc_if_i[22] ),
    .QN(_13531_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(_01389_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_if_i[23] ),
    .QN(_13530_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(_01390_),
    .CK(clknet_leaf_43_clk),
    .Q(\cs_registers_i.pc_if_i[24] ),
    .QN(_13529_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(_01391_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[25] ),
    .QN(_13528_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(_01392_),
    .CK(clknet_leaf_43_clk),
    .Q(\cs_registers_i.pc_if_i[26] ),
    .QN(_13527_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(_01393_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[27] ),
    .QN(_13526_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(_01394_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[28] ),
    .QN(_13525_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(_01395_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[29] ),
    .QN(_13524_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(_01396_),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.pc_if_i[30] ),
    .QN(_13523_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(_01397_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[3] ),
    .QN(_13522_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(_01398_),
    .CK(clknet_leaf_47_clk),
    .Q(\cs_registers_i.pc_if_i[31] ),
    .QN(_13521_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(_01399_),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.pc_if_i[4] ),
    .QN(_13520_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(_01400_),
    .CK(clknet_leaf_46_clk),
    .Q(\cs_registers_i.pc_if_i[5] ),
    .QN(_13519_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(_01401_),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.pc_if_i[6] ),
    .QN(_13518_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(_01402_),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.pc_if_i[7] ),
    .QN(_13517_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(_01403_),
    .CK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.pc_if_i[8] ),
    .QN(_13516_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(_01404_),
    .CK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.pc_if_i[9] ),
    .QN(_13515_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(_01405_),
    .CK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.pc_if_i[10] ),
    .QN(_13514_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(_01406_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .QN(_13513_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(_01407_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .QN(_13512_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(_01408_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .QN(_13511_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(_01409_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .QN(_13510_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(_01410_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .QN(_13509_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(_01411_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .QN(_13508_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(_01412_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .QN(_13507_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(_01413_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .QN(_13506_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(_01414_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .QN(_13505_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(_01415_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .QN(_13504_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(_01416_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .QN(_13503_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(_01417_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .QN(_13502_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(_01418_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .QN(_13501_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(_01419_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .QN(_13500_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(_01420_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .QN(_13499_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(_01421_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .QN(_13498_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(_01422_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .QN(_13497_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(_01423_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .QN(_13496_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(_01424_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .QN(_13495_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(_01425_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .QN(_13494_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(_01426_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .QN(_13493_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(_01427_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .QN(_13492_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(_01428_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .QN(_13491_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(_01429_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .QN(_13490_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(_01430_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .QN(_13489_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(_01431_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .QN(_13488_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(_01432_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .QN(_13487_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(_01433_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .QN(_13486_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(_01434_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .QN(_13485_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(_01435_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .QN(_13484_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(_01436_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .QN(_13483_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(_01437_),
    .CK(clknet_leaf_127_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .QN(_13482_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(_01438_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .QN(_13481_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(_01439_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .QN(_13480_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(_01440_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .QN(_13479_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(_01441_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .QN(_13478_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(_01442_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .QN(_13477_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(_01443_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .QN(_13476_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(_01444_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .QN(_13475_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(_01445_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .QN(_13474_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(_01446_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .QN(_13473_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(_01447_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .QN(_13472_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(_01448_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .QN(_13471_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(_01449_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .QN(_13470_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(_01450_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .QN(_13469_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(_01451_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .QN(_13468_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(_01452_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .QN(_13467_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(_01453_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .QN(_13466_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(_01454_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .QN(_13465_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(_01455_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .QN(_13464_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(_01456_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .QN(_13463_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(_01457_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .QN(_13462_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(_01458_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .QN(_13461_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(_01459_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .QN(_13460_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(_01460_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .QN(_13459_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(_01461_),
    .CK(clknet_leaf_127_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .QN(_13458_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(_01462_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .QN(_13457_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(_01463_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .QN(_13456_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(_01464_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .QN(_13455_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(_01465_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .QN(_13454_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(_01466_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .QN(_13453_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(_01467_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .QN(_13452_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(_01468_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .QN(_13451_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(_01469_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .QN(_13450_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(_01470_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .QN(_13449_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(_01471_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .QN(_13448_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(_01472_),
    .CK(clknet_leaf_127_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .QN(_13447_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(_01473_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .QN(_13446_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(_01474_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .QN(_13445_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(_01475_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .QN(_13444_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(_01476_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .QN(_13443_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(_01477_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .QN(_13442_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(_01478_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .QN(_13441_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(_01479_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .QN(_13440_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(_01480_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .QN(_13439_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(_01481_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .QN(_13438_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(_01482_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .QN(_13437_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(_01483_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .QN(_13436_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(_01484_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .QN(_13435_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(_01485_),
    .CK(clknet_leaf_134_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .QN(_13434_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(_01486_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .QN(_13433_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(_01487_),
    .CK(clknet_leaf_130_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .QN(_13432_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(_01488_),
    .CK(clknet_leaf_129_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .QN(_13431_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(_01489_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .QN(_13430_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(_01490_),
    .CK(clknet_leaf_128_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .QN(_13429_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(_01491_),
    .CK(clknet_leaf_123_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .QN(_13428_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(_01492_),
    .CK(clknet_leaf_124_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .QN(_13427_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(_01493_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .QN(_13426_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(_01494_),
    .CK(clknet_leaf_125_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .QN(_13425_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(_01495_),
    .CK(clknet_leaf_133_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .QN(_13424_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(_01496_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .QN(_13423_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(_01497_),
    .CK(clknet_leaf_132_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .QN(_13422_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(_01498_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .QN(_13421_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(_01499_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .QN(_13420_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(_01500_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .QN(_13419_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(_01501_),
    .CK(clknet_leaf_131_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .QN(_14060_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .RN(net261),
    .CK(clknet_leaf_126_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .QN(_00136_));
 DFFR_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .RN(net261),
    .CK(clknet_leaf_115_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .QN(_00135_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .RN(net261),
    .CK(clknet_leaf_115_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .QN(_14061_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .RN(net261),
    .CK(clknet_leaf_111_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .QN(_14062_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .RN(net261),
    .CK(clknet_leaf_111_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .QN(_00134_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(_01502_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .QN(_13418_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(_01503_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .QN(_13417_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(_01504_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .QN(_13416_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(_01505_),
    .CK(clknet_leaf_40_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .QN(_13415_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(_01506_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .QN(_13414_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(_01507_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .QN(_13413_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(_01508_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .QN(_13412_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(_01509_),
    .CK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .QN(_13411_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(_01510_),
    .CK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .QN(_13410_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(_01511_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .QN(_13409_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(_01512_),
    .CK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .QN(_13408_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(_01513_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .QN(_13407_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(_01514_),
    .CK(clknet_leaf_33_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .QN(_13406_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(_01515_),
    .CK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .QN(_13405_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(_01516_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .QN(_13404_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(_01517_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .QN(_13403_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(_01518_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .QN(_13402_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(_01519_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .QN(_13401_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(_01520_),
    .CK(clknet_leaf_33_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .QN(_13400_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(_01521_),
    .CK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .QN(_13399_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(_01522_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .QN(_13398_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(_01523_),
    .CK(clknet_leaf_34_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .QN(_13397_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(_01524_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .QN(_13396_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(_01525_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .QN(_13395_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(_01526_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .QN(_13394_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(_01527_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .QN(_13393_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(_01528_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .QN(_13392_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(_01529_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .QN(_13391_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(_01530_),
    .CK(clknet_leaf_42_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .QN(_13390_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(_01531_),
    .CK(clknet_leaf_41_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .QN(_14063_));
 DFFR_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .RN(net261),
    .CK(clknet_leaf_110_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .QN(_00133_));
 DFF_X1 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(_01532_),
    .CK(clknet_leaf_127_clk),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .QN(_13389_));
 DFF_X1 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(_01533_),
    .CK(clknet_leaf_111_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ),
    .QN(_13388_));
 DFF_X1 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_01534_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .QN(_13387_));
 DFF_X1 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(_01535_),
    .CK(clknet_leaf_6_clk),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ),
    .QN(_00278_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[0]$_DFFE_PN_  (.D(_01536_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_i[0] ),
    .QN(_13386_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[10]$_DFFE_PN_  (.D(_01537_),
    .CK(clknet_leaf_8_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .QN(_00036_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[11]$_DFFE_PN_  (.D(_01538_),
    .CK(clknet_leaf_6_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .QN(_00039_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[12]$_DFFE_PN_  (.D(_01539_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_i[12] ),
    .QN(_00176_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[13]$_DFFE_PN_  (.D(_01540_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_i[13] ),
    .QN(_00175_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[14]$_DFFE_PN_  (.D(_01541_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_i[14] ),
    .QN(_00173_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[15]$_DFFE_PN_  (.D(_01542_),
    .CK(clknet_leaf_5_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .QN(_00184_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[16]$_DFFE_PN_  (.D(_01543_),
    .CK(clknet_leaf_5_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .QN(_00183_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[17]$_DFFE_PN_  (.D(_01544_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .QN(_00182_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[18]$_DFFE_PN_  (.D(_01545_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .QN(_00181_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[19]$_DFFE_PN_  (.D(_01546_),
    .CK(clknet_leaf_5_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .QN(_00180_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[1]$_DFFE_PN_  (.D(_01547_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[1] ),
    .QN(_00013_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[20]$_DFFE_PN_  (.D(_01548_),
    .CK(clknet_leaf_6_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .QN(_00140_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[21]$_DFFE_PN_  (.D(_01549_),
    .CK(clknet_leaf_11_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .QN(_13385_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[22]$_DFFE_PN_  (.D(_01550_),
    .CK(clknet_leaf_5_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .QN(_13384_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[23]$_DFFE_PN_  (.D(_01551_),
    .CK(clknet_leaf_5_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .QN(_00139_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[24]$_DFFE_PN_  (.D(_01552_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .QN(_00138_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[25]$_DFFE_PN_  (.D(_01553_),
    .CK(clknet_leaf_5_clk),
    .Q(\id_stage_i.controller_i.instr_i[25] ),
    .QN(_13383_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[26]$_DFFE_PN_  (.D(_01554_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_i[26] ),
    .QN(_00177_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[27]$_DFFE_PN_  (.D(_01555_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[27] ),
    .QN(_13382_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[28]$_DFFE_PN_  (.D(_01556_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[28] ),
    .QN(_13381_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[29]$_DFFE_PN_  (.D(_01557_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[29] ),
    .QN(_13380_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[2]$_DFFE_PN_  (.D(_01558_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_i[2] ),
    .QN(_00015_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[30]$_DFFE_PN_  (.D(_01559_),
    .CK(clknet_leaf_5_clk),
    .Q(\id_stage_i.controller_i.instr_i[30] ),
    .QN(_13379_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[31]$_DFFE_PN_  (.D(_01560_),
    .CK(clknet_leaf_5_clk),
    .Q(\id_stage_i.controller_i.instr_i[31] ),
    .QN(_00174_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[3]$_DFFE_PN_  (.D(_01561_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_i[3] ),
    .QN(_00017_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[4]$_DFFE_PN_  (.D(_01562_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_i[4] ),
    .QN(_00020_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[5]$_DFFE_PN_  (.D(_01563_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_i[5] ),
    .QN(_00023_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[6]$_DFFE_PN_  (.D(_01564_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_i[6] ),
    .QN(_00172_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[7]$_DFFE_PN_  (.D(_01565_),
    .CK(clknet_leaf_9_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .QN(_00216_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[8]$_DFFE_PN_  (.D(_01566_),
    .CK(clknet_leaf_8_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .QN(_00030_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[9]$_DFFE_PN_  (.D(_01567_),
    .CK(clknet_leaf_8_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .QN(_00033_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(_01568_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .QN(_13378_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(_01569_),
    .CK(clknet_leaf_127_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .QN(_00037_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_01570_),
    .CK(clknet_leaf_2_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .QN(_00040_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_01571_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .QN(_00042_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_01572_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .QN(_00044_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_01573_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .QN(_00046_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_01574_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .QN(_00048_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_01575_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .QN(_00014_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(_01576_),
    .CK(clknet_leaf_113_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .QN(_00016_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(_01577_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .QN(_00018_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(_01578_),
    .CK(clknet_leaf_115_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .QN(_00021_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(_01579_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .QN(_00024_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(_01580_),
    .CK(clknet_leaf_115_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .QN(_00026_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(_01581_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .QN(_00028_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_01582_),
    .CK(clknet_leaf_114_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .QN(_00031_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(_01583_),
    .CK(clknet_leaf_112_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .QN(_00034_));
 DFFR_X2 \if_stage_i.instr_valid_id_q$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .RN(net262),
    .CK(clknet_leaf_110_clk),
    .Q(\id_stage_i.controller_i.instr_valid_i ),
    .QN(_01161_));
 DFF_X1 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(_01584_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[10] ),
    .QN(_00038_));
 DFF_X1 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(_01585_),
    .CK(clknet_leaf_54_clk),
    .Q(\cs_registers_i.pc_id_i[11] ),
    .QN(_00041_));
 DFF_X2 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(_01586_),
    .CK(clknet_leaf_54_clk),
    .Q(\cs_registers_i.pc_id_i[12] ),
    .QN(_00043_));
 DFF_X1 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(_01587_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[13] ),
    .QN(_00045_));
 DFF_X1 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(_01588_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[14] ),
    .QN(_00047_));
 DFF_X1 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(_01589_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[15] ),
    .QN(_00049_));
 DFF_X1 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(_01590_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[16] ),
    .QN(_00050_));
 DFF_X2 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(_01591_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[17] ),
    .QN(_00051_));
 DFF_X2 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(_01592_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[18] ),
    .QN(_00052_));
 DFF_X1 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(_01593_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[19] ),
    .QN(_00053_));
 DFF_X1 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(_01594_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[1] ),
    .QN(_13377_));
 DFF_X1 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(_01595_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[20] ),
    .QN(_00054_));
 DFF_X2 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(_01596_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[21] ),
    .QN(_00055_));
 DFF_X2 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(_01597_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[22] ),
    .QN(_00056_));
 DFF_X1 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(_01598_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[23] ),
    .QN(_00057_));
 DFF_X1 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(_01599_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[24] ),
    .QN(_00058_));
 DFF_X1 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(_01600_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[25] ),
    .QN(_00059_));
 DFF_X1 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(_01601_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_id_i[26] ),
    .QN(_00060_));
 DFF_X1 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(_01602_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_id_i[27] ),
    .QN(_00061_));
 DFF_X2 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(_01603_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_id_i[28] ),
    .QN(_00062_));
 DFF_X2 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(_01604_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_id_i[29] ),
    .QN(_00063_));
 DFF_X2 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(_01605_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_id_i[2] ),
    .QN(_00012_));
 DFF_X1 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(_01606_),
    .CK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.pc_id_i[30] ),
    .QN(_00064_));
 DFF_X1 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(_01607_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_id_i[31] ),
    .QN(_00065_));
 DFF_X1 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(_01608_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[3] ),
    .QN(_00019_));
 DFF_X1 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(_01609_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[4] ),
    .QN(_00022_));
 DFF_X1 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(_01610_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[5] ),
    .QN(_00025_));
 DFF_X1 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(_01611_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[6] ),
    .QN(_00027_));
 DFF_X1 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(_01612_),
    .CK(clknet_leaf_55_clk),
    .Q(\cs_registers_i.pc_id_i[7] ),
    .QN(_00029_));
 DFF_X1 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(_01613_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[8] ),
    .QN(_00032_));
 DFF_X1 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(_01614_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[9] ),
    .QN(_00035_));
 DFFR_X2 \load_store_unit_i.addr_last_q[0]$_DFFE_PN0P_  (.D(_01615_),
    .RN(net264),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .QN(_13376_));
 DFFR_X1 \load_store_unit_i.addr_last_q[10]$_DFFE_PN0P_  (.D(_01616_),
    .RN(net264),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .QN(_13375_));
 DFFR_X1 \load_store_unit_i.addr_last_q[11]$_DFFE_PN0P_  (.D(_01617_),
    .RN(net264),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .QN(_13374_));
 DFFR_X1 \load_store_unit_i.addr_last_q[12]$_DFFE_PN0P_  (.D(_01618_),
    .RN(net264),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .QN(_13373_));
 DFFR_X2 \load_store_unit_i.addr_last_q[13]$_DFFE_PN0P_  (.D(_01619_),
    .RN(net264),
    .CK(clknet_leaf_22_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .QN(_13372_));
 DFFR_X2 \load_store_unit_i.addr_last_q[14]$_DFFE_PN0P_  (.D(_01620_),
    .RN(net264),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .QN(_13371_));
 DFFR_X2 \load_store_unit_i.addr_last_q[15]$_DFFE_PN0P_  (.D(_01621_),
    .RN(net264),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .QN(_13370_));
 DFFR_X1 \load_store_unit_i.addr_last_q[16]$_DFFE_PN0P_  (.D(_01622_),
    .RN(net264),
    .CK(clknet_leaf_22_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .QN(_13369_));
 DFFR_X1 \load_store_unit_i.addr_last_q[17]$_DFFE_PN0P_  (.D(_01623_),
    .RN(net264),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .QN(_13368_));
 DFFR_X2 \load_store_unit_i.addr_last_q[18]$_DFFE_PN0P_  (.D(_01624_),
    .RN(net264),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .QN(_13367_));
 DFFR_X1 \load_store_unit_i.addr_last_q[19]$_DFFE_PN0P_  (.D(_01625_),
    .RN(net264),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .QN(_13366_));
 DFFR_X2 \load_store_unit_i.addr_last_q[1]$_DFFE_PN0P_  (.D(_01626_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .QN(_13365_));
 DFFR_X2 \load_store_unit_i.addr_last_q[20]$_DFFE_PN0P_  (.D(_01627_),
    .RN(net264),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .QN(_13364_));
 DFFR_X2 \load_store_unit_i.addr_last_q[21]$_DFFE_PN0P_  (.D(_01628_),
    .RN(net264),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .QN(_13363_));
 DFFR_X1 \load_store_unit_i.addr_last_q[22]$_DFFE_PN0P_  (.D(_01629_),
    .RN(net264),
    .CK(clknet_leaf_22_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .QN(_13362_));
 DFFR_X1 \load_store_unit_i.addr_last_q[23]$_DFFE_PN0P_  (.D(_01630_),
    .RN(net264),
    .CK(clknet_leaf_22_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .QN(_13361_));
 DFFR_X1 \load_store_unit_i.addr_last_q[24]$_DFFE_PN0P_  (.D(_01631_),
    .RN(net264),
    .CK(clknet_leaf_22_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .QN(_13360_));
 DFFR_X1 \load_store_unit_i.addr_last_q[25]$_DFFE_PN0P_  (.D(_01632_),
    .RN(net264),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .QN(_13359_));
 DFFR_X1 \load_store_unit_i.addr_last_q[26]$_DFFE_PN0P_  (.D(_01633_),
    .RN(net264),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .QN(_13358_));
 DFFR_X2 \load_store_unit_i.addr_last_q[27]$_DFFE_PN0P_  (.D(_01634_),
    .RN(net264),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .QN(_13357_));
 DFFR_X1 \load_store_unit_i.addr_last_q[28]$_DFFE_PN0P_  (.D(_01635_),
    .RN(net264),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .QN(_13356_));
 DFFR_X1 \load_store_unit_i.addr_last_q[29]$_DFFE_PN0P_  (.D(_01636_),
    .RN(net264),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .QN(_13355_));
 DFFR_X1 \load_store_unit_i.addr_last_q[2]$_DFFE_PN0P_  (.D(_01637_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .QN(_13354_));
 DFFR_X1 \load_store_unit_i.addr_last_q[30]$_DFFE_PN0P_  (.D(_01638_),
    .RN(net264),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .QN(_13353_));
 DFFR_X1 \load_store_unit_i.addr_last_q[31]$_DFFE_PN0P_  (.D(_01639_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .QN(_13352_));
 DFFR_X1 \load_store_unit_i.addr_last_q[3]$_DFFE_PN0P_  (.D(_01640_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .QN(_13351_));
 DFFR_X1 \load_store_unit_i.addr_last_q[4]$_DFFE_PN0P_  (.D(_01641_),
    .RN(net264),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .QN(_13350_));
 DFFR_X2 \load_store_unit_i.addr_last_q[5]$_DFFE_PN0P_  (.D(_01642_),
    .RN(net264),
    .CK(clknet_leaf_58_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .QN(_13349_));
 DFFR_X1 \load_store_unit_i.addr_last_q[6]$_DFFE_PN0P_  (.D(_01643_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .QN(_13348_));
 DFFR_X1 \load_store_unit_i.addr_last_q[7]$_DFFE_PN0P_  (.D(_01644_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .QN(_13347_));
 DFFR_X1 \load_store_unit_i.addr_last_q[8]$_DFFE_PN0P_  (.D(_01645_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .QN(_13346_));
 DFFR_X1 \load_store_unit_i.addr_last_q[9]$_DFFE_PN0P_  (.D(_01646_),
    .RN(net264),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .QN(_13345_));
 DFFR_X2 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_01647_),
    .RN(net260),
    .CK(clknet_leaf_9_clk),
    .Q(\load_store_unit_i.data_sign_ext_q ),
    .QN(_13344_));
 DFFR_X2 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_01648_),
    .RN(net260),
    .CK(clknet_leaf_9_clk),
    .Q(\load_store_unit_i.data_we_q ),
    .QN(_01160_));
 DFFR_X2 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_01649_),
    .RN(net260),
    .CK(clknet_leaf_6_clk),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .QN(_16085_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_01650_),
    .RN(net260),
    .CK(clknet_leaf_6_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ),
    .QN(_13343_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_01651_),
    .RN(net260),
    .CK(clknet_leaf_6_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ),
    .QN(_13342_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_01652_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ),
    .QN(_00171_));
 DFFR_X1 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_01653_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.lsu_err_q ),
    .QN(_13341_));
 DFFR_X1 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_01654_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.rdata_offset_q[0] ),
    .QN(_13340_));
 DFFR_X1 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_01655_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.rdata_offset_q[1] ),
    .QN(_13339_));
 DFFR_X1 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_01656_),
    .RN(net255),
    .CK(clknet_leaf_1_clk),
    .Q(\load_store_unit_i.rdata_q[8] ),
    .QN(_13338_));
 DFFR_X1 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_01657_),
    .RN(net255),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[18] ),
    .QN(_13337_));
 DFFR_X1 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_01658_),
    .RN(net255),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[19] ),
    .QN(_13336_));
 DFFR_X1 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_01659_),
    .RN(net255),
    .CK(clknet_leaf_0_clk),
    .Q(\load_store_unit_i.rdata_q[20] ),
    .QN(_13335_));
 DFFR_X1 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_01660_),
    .RN(net255),
    .CK(clknet_leaf_0_clk),
    .Q(\load_store_unit_i.rdata_q[21] ),
    .QN(_13334_));
 DFFR_X1 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_01661_),
    .RN(net260),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[22] ),
    .QN(_13333_));
 DFFR_X1 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_01662_),
    .RN(net261),
    .CK(clknet_leaf_2_clk),
    .Q(\load_store_unit_i.rdata_q[23] ),
    .QN(_13332_));
 DFFR_X1 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_01663_),
    .RN(net255),
    .CK(clknet_leaf_2_clk),
    .Q(\load_store_unit_i.rdata_q[24] ),
    .QN(_13331_));
 DFFR_X1 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_01664_),
    .RN(net260),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[25] ),
    .QN(_13330_));
 DFFR_X1 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_01665_),
    .RN(net260),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[26] ),
    .QN(_13329_));
 DFFR_X1 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_01666_),
    .RN(net255),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[27] ),
    .QN(_13328_));
 DFFR_X1 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_01667_),
    .RN(net260),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[9] ),
    .QN(_13327_));
 DFFR_X1 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_01668_),
    .RN(net255),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[28] ),
    .QN(_13326_));
 DFFR_X1 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_01669_),
    .RN(net255),
    .CK(clknet_leaf_1_clk),
    .Q(\load_store_unit_i.rdata_q[29] ),
    .QN(_13325_));
 DFFR_X1 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_01670_),
    .RN(net260),
    .CK(clknet_leaf_7_clk),
    .Q(\load_store_unit_i.rdata_q[30] ),
    .QN(_13324_));
 DFFR_X1 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_01671_),
    .RN(net260),
    .CK(clknet_leaf_8_clk),
    .Q(\load_store_unit_i.rdata_q[31] ),
    .QN(_13323_));
 DFFR_X1 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_01672_),
    .RN(net255),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[10] ),
    .QN(_13322_));
 DFFR_X1 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_01673_),
    .RN(net255),
    .CK(clknet_leaf_4_clk),
    .Q(\load_store_unit_i.rdata_q[11] ),
    .QN(_13321_));
 DFFR_X1 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_01674_),
    .RN(net255),
    .CK(clknet_leaf_0_clk),
    .Q(\load_store_unit_i.rdata_q[12] ),
    .QN(_13320_));
 DFFR_X1 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_01675_),
    .RN(net255),
    .CK(clknet_leaf_1_clk),
    .Q(\load_store_unit_i.rdata_q[13] ),
    .QN(_13319_));
 DFFR_X1 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_01676_),
    .RN(net260),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[14] ),
    .QN(_13318_));
 DFFR_X1 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_01677_),
    .RN(net261),
    .CK(clknet_leaf_2_clk),
    .Q(\load_store_unit_i.rdata_q[15] ),
    .QN(_13317_));
 DFFR_X1 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_01678_),
    .RN(net255),
    .CK(clknet_leaf_2_clk),
    .Q(\load_store_unit_i.rdata_q[16] ),
    .QN(_13316_));
 DFFR_X1 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_01679_),
    .RN(net260),
    .CK(clknet_leaf_3_clk),
    .Q(\load_store_unit_i.rdata_q[17] ),
    .QN(_13315_));
 NOR2_X4 clone1 (.A1(_03792_),
    .A2(_03662_),
    .ZN(net1));
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_425 ();
 BUF_X4 max_cap12 (.A(\alu_adder_result_ex[29] ),
    .Z(net14));
 BUF_X8 max_cap13 (.A(\alu_adder_result_ex[1] ),
    .Z(net15));
 BUF_X4 max_cap14 (.A(_04510_),
    .Z(net16));
 BUF_X4 max_cap15 (.A(_05198_),
    .Z(net17));
 BUF_X2 max_cap16 (.A(net19),
    .Z(net18));
 BUF_X4 max_cap17 (.A(net20),
    .Z(net19));
 CLKBUF_X3 wire18 (.A(_10391_),
    .Z(net20));
 CLKBUF_X2 wire19 (.A(_11489_),
    .Z(net21));
 BUF_X4 max_cap20 (.A(_03437_),
    .Z(net22));
 BUF_X1 input1 (.A(boot_addr_i[10]),
    .Z(net3));
 BUF_X1 input2 (.A(boot_addr_i[11]),
    .Z(net4));
 CLKBUF_X2 input3 (.A(boot_addr_i[12]),
    .Z(net5));
 BUF_X1 input4 (.A(boot_addr_i[13]),
    .Z(net6));
 BUF_X1 input5 (.A(boot_addr_i[14]),
    .Z(net7));
 CLKBUF_X2 input6 (.A(boot_addr_i[15]),
    .Z(net8));
 BUF_X1 input7 (.A(boot_addr_i[16]),
    .Z(net9));
 CLKBUF_X2 input8 (.A(boot_addr_i[17]),
    .Z(net10));
 BUF_X2 input9 (.A(boot_addr_i[18]),
    .Z(net11));
 BUF_X1 input10 (.A(boot_addr_i[19]),
    .Z(net12));
 BUF_X1 input11 (.A(boot_addr_i[20]),
    .Z(net13));
 BUF_X1 input12 (.A(boot_addr_i[21]),
    .Z(net23));
 BUF_X1 input13 (.A(boot_addr_i[22]),
    .Z(net24));
 CLKBUF_X2 input14 (.A(boot_addr_i[23]),
    .Z(net25));
 BUF_X1 input15 (.A(boot_addr_i[24]),
    .Z(net26));
 BUF_X1 input16 (.A(boot_addr_i[25]),
    .Z(net27));
 BUF_X1 input17 (.A(boot_addr_i[26]),
    .Z(net28));
 BUF_X1 input18 (.A(boot_addr_i[27]),
    .Z(net29));
 BUF_X1 input19 (.A(boot_addr_i[28]),
    .Z(net30));
 BUF_X1 input20 (.A(boot_addr_i[29]),
    .Z(net31));
 BUF_X1 input21 (.A(boot_addr_i[30]),
    .Z(net32));
 CLKBUF_X2 input22 (.A(boot_addr_i[31]),
    .Z(net33));
 BUF_X1 input23 (.A(boot_addr_i[8]),
    .Z(net34));
 BUF_X1 input24 (.A(boot_addr_i[9]),
    .Z(net35));
 BUF_X2 input25 (.A(data_err_i),
    .Z(net36));
 CLKBUF_X3 input26 (.A(data_gnt_i),
    .Z(net37));
 BUF_X2 input27 (.A(data_rdata_i[0]),
    .Z(net38));
 BUF_X2 input28 (.A(data_rdata_i[10]),
    .Z(net39));
 BUF_X2 input29 (.A(data_rdata_i[11]),
    .Z(net40));
 CLKBUF_X2 input30 (.A(data_rdata_i[12]),
    .Z(net41));
 CLKBUF_X2 input31 (.A(data_rdata_i[13]),
    .Z(net42));
 BUF_X2 input32 (.A(data_rdata_i[14]),
    .Z(net43));
 BUF_X2 input33 (.A(data_rdata_i[15]),
    .Z(net44));
 BUF_X1 input34 (.A(data_rdata_i[16]),
    .Z(net45));
 BUF_X2 input35 (.A(data_rdata_i[17]),
    .Z(net46));
 BUF_X2 input36 (.A(data_rdata_i[18]),
    .Z(net47));
 BUF_X2 input37 (.A(data_rdata_i[19]),
    .Z(net48));
 BUF_X2 input38 (.A(data_rdata_i[1]),
    .Z(net49));
 CLKBUF_X2 input39 (.A(data_rdata_i[20]),
    .Z(net50));
 CLKBUF_X2 input40 (.A(data_rdata_i[21]),
    .Z(net51));
 BUF_X2 input41 (.A(data_rdata_i[22]),
    .Z(net52));
 CLKBUF_X2 input42 (.A(data_rdata_i[24]),
    .Z(net53));
 BUF_X2 input43 (.A(data_rdata_i[25]),
    .Z(net54));
 BUF_X2 input44 (.A(data_rdata_i[26]),
    .Z(net55));
 BUF_X2 input45 (.A(data_rdata_i[27]),
    .Z(net56));
 CLKBUF_X2 input46 (.A(data_rdata_i[28]),
    .Z(net57));
 CLKBUF_X2 input47 (.A(data_rdata_i[29]),
    .Z(net58));
 BUF_X2 input48 (.A(data_rdata_i[2]),
    .Z(net59));
 BUF_X2 input49 (.A(data_rdata_i[30]),
    .Z(net60));
 BUF_X2 input50 (.A(data_rdata_i[31]),
    .Z(net61));
 BUF_X2 input51 (.A(data_rdata_i[3]),
    .Z(net62));
 BUF_X1 input52 (.A(data_rdata_i[4]),
    .Z(net63));
 BUF_X1 input53 (.A(data_rdata_i[5]),
    .Z(net64));
 BUF_X2 input54 (.A(data_rdata_i[6]),
    .Z(net65));
 BUF_X2 input55 (.A(data_rdata_i[7]),
    .Z(net66));
 BUF_X2 input56 (.A(data_rdata_i[8]),
    .Z(net67));
 BUF_X2 input57 (.A(data_rdata_i[9]),
    .Z(net68));
 BUF_X2 input58 (.A(debug_req_i),
    .Z(net69));
 BUF_X1 input59 (.A(fetch_enable_i),
    .Z(net70));
 BUF_X1 input60 (.A(hart_id_i[0]),
    .Z(net71));
 BUF_X1 input61 (.A(hart_id_i[10]),
    .Z(net72));
 BUF_X1 input62 (.A(hart_id_i[11]),
    .Z(net73));
 BUF_X1 input63 (.A(hart_id_i[12]),
    .Z(net74));
 BUF_X1 input64 (.A(hart_id_i[13]),
    .Z(net75));
 BUF_X1 input65 (.A(hart_id_i[14]),
    .Z(net76));
 BUF_X1 input66 (.A(hart_id_i[15]),
    .Z(net77));
 BUF_X1 input67 (.A(hart_id_i[16]),
    .Z(net78));
 BUF_X1 input68 (.A(hart_id_i[17]),
    .Z(net79));
 BUF_X1 input69 (.A(hart_id_i[18]),
    .Z(net80));
 BUF_X1 input70 (.A(hart_id_i[19]),
    .Z(net81));
 BUF_X1 input71 (.A(hart_id_i[1]),
    .Z(net82));
 BUF_X1 input72 (.A(hart_id_i[20]),
    .Z(net83));
 BUF_X1 input73 (.A(hart_id_i[21]),
    .Z(net84));
 BUF_X1 input74 (.A(hart_id_i[22]),
    .Z(net85));
 BUF_X1 input75 (.A(hart_id_i[23]),
    .Z(net86));
 BUF_X1 input76 (.A(hart_id_i[24]),
    .Z(net87));
 BUF_X1 input77 (.A(hart_id_i[25]),
    .Z(net88));
 BUF_X1 input78 (.A(hart_id_i[26]),
    .Z(net89));
 BUF_X1 input79 (.A(hart_id_i[27]),
    .Z(net90));
 BUF_X1 input80 (.A(hart_id_i[28]),
    .Z(net91));
 BUF_X1 input81 (.A(hart_id_i[29]),
    .Z(net92));
 BUF_X1 input82 (.A(hart_id_i[2]),
    .Z(net93));
 BUF_X1 input83 (.A(hart_id_i[30]),
    .Z(net94));
 BUF_X1 input84 (.A(hart_id_i[31]),
    .Z(net95));
 BUF_X1 input85 (.A(hart_id_i[3]),
    .Z(net96));
 BUF_X1 input86 (.A(hart_id_i[4]),
    .Z(net97));
 BUF_X1 input87 (.A(hart_id_i[5]),
    .Z(net98));
 BUF_X1 input88 (.A(hart_id_i[6]),
    .Z(net99));
 BUF_X1 input89 (.A(hart_id_i[7]),
    .Z(net100));
 BUF_X1 input90 (.A(hart_id_i[8]),
    .Z(net101));
 BUF_X1 input91 (.A(hart_id_i[9]),
    .Z(net102));
 CLKBUF_X3 input92 (.A(instr_gnt_i),
    .Z(net103));
 BUF_X1 input93 (.A(instr_rdata_i[0]),
    .Z(net104));
 BUF_X1 input94 (.A(instr_rdata_i[10]),
    .Z(net105));
 BUF_X1 input95 (.A(instr_rdata_i[11]),
    .Z(net106));
 BUF_X1 input96 (.A(instr_rdata_i[12]),
    .Z(net107));
 BUF_X1 input97 (.A(instr_rdata_i[13]),
    .Z(net108));
 BUF_X1 input98 (.A(instr_rdata_i[14]),
    .Z(net109));
 BUF_X1 input99 (.A(instr_rdata_i[15]),
    .Z(net110));
 BUF_X1 input100 (.A(instr_rdata_i[18]),
    .Z(net111));
 BUF_X1 input101 (.A(instr_rdata_i[19]),
    .Z(net112));
 BUF_X1 input102 (.A(instr_rdata_i[1]),
    .Z(net113));
 BUF_X1 input103 (.A(instr_rdata_i[20]),
    .Z(net114));
 BUF_X1 input104 (.A(instr_rdata_i[21]),
    .Z(net115));
 BUF_X1 input105 (.A(instr_rdata_i[22]),
    .Z(net116));
 BUF_X1 input106 (.A(instr_rdata_i[23]),
    .Z(net117));
 BUF_X1 input107 (.A(instr_rdata_i[24]),
    .Z(net118));
 BUF_X1 input108 (.A(instr_rdata_i[25]),
    .Z(net119));
 BUF_X1 input109 (.A(instr_rdata_i[26]),
    .Z(net120));
 BUF_X1 input110 (.A(instr_rdata_i[27]),
    .Z(net121));
 BUF_X1 input111 (.A(instr_rdata_i[28]),
    .Z(net122));
 BUF_X1 input112 (.A(instr_rdata_i[29]),
    .Z(net123));
 BUF_X1 input113 (.A(instr_rdata_i[2]),
    .Z(net124));
 CLKBUF_X2 input114 (.A(instr_rdata_i[30]),
    .Z(net125));
 CLKBUF_X2 input115 (.A(instr_rdata_i[31]),
    .Z(net126));
 BUF_X1 input116 (.A(instr_rdata_i[3]),
    .Z(net127));
 BUF_X1 input117 (.A(instr_rdata_i[4]),
    .Z(net128));
 BUF_X1 input118 (.A(instr_rdata_i[5]),
    .Z(net129));
 BUF_X1 input119 (.A(instr_rdata_i[6]),
    .Z(net130));
 BUF_X1 input120 (.A(instr_rdata_i[7]),
    .Z(net131));
 BUF_X1 input121 (.A(instr_rdata_i[8]),
    .Z(net132));
 BUF_X1 input122 (.A(instr_rdata_i[9]),
    .Z(net133));
 CLKBUF_X2 input123 (.A(instr_rvalid_i),
    .Z(net134));
 BUF_X2 input124 (.A(irq_external_i),
    .Z(net135));
 BUF_X2 input125 (.A(irq_fast_i[0]),
    .Z(net136));
 BUF_X1 input126 (.A(irq_fast_i[10]),
    .Z(net137));
 BUF_X1 input127 (.A(irq_fast_i[11]),
    .Z(net138));
 BUF_X2 input128 (.A(irq_fast_i[12]),
    .Z(net139));
 BUF_X2 input129 (.A(irq_fast_i[13]),
    .Z(net140));
 BUF_X1 input130 (.A(irq_fast_i[14]),
    .Z(net141));
 BUF_X2 input131 (.A(irq_fast_i[1]),
    .Z(net142));
 BUF_X2 input132 (.A(irq_fast_i[2]),
    .Z(net143));
 BUF_X2 input133 (.A(irq_fast_i[3]),
    .Z(net144));
 BUF_X2 input134 (.A(irq_fast_i[4]),
    .Z(net145));
 CLKBUF_X2 input135 (.A(irq_fast_i[5]),
    .Z(net146));
 BUF_X2 input136 (.A(irq_fast_i[6]),
    .Z(net147));
 BUF_X2 input137 (.A(irq_fast_i[7]),
    .Z(net148));
 BUF_X1 input138 (.A(irq_fast_i[8]),
    .Z(net149));
 CLKBUF_X2 input139 (.A(irq_fast_i[9]),
    .Z(net150));
 BUF_X2 input140 (.A(irq_software_i),
    .Z(net151));
 BUF_X1 input141 (.A(irq_timer_i),
    .Z(net152));
 BUF_X32 input142 (.A(net387),
    .Z(net153));
 BUF_X1 input143 (.A(test_en_i),
    .Z(net154));
 BUF_X1 output144 (.A(net155),
    .Z(core_sleep_o));
 BUF_X1 output145 (.A(net156),
    .Z(data_addr_o[10]));
 BUF_X1 output146 (.A(net157),
    .Z(data_addr_o[11]));
 BUF_X1 output147 (.A(net158),
    .Z(data_addr_o[12]));
 BUF_X1 output148 (.A(net159),
    .Z(data_addr_o[13]));
 BUF_X1 output149 (.A(net160),
    .Z(data_addr_o[14]));
 BUF_X1 output150 (.A(net161),
    .Z(data_addr_o[15]));
 BUF_X1 output151 (.A(net162),
    .Z(data_addr_o[16]));
 BUF_X1 output152 (.A(net163),
    .Z(data_addr_o[17]));
 BUF_X1 output153 (.A(net164),
    .Z(data_addr_o[18]));
 BUF_X1 output154 (.A(net165),
    .Z(data_addr_o[19]));
 BUF_X1 output155 (.A(net166),
    .Z(data_addr_o[20]));
 BUF_X1 output156 (.A(net167),
    .Z(data_addr_o[21]));
 BUF_X1 output157 (.A(net168),
    .Z(data_addr_o[22]));
 BUF_X1 output158 (.A(net169),
    .Z(data_addr_o[23]));
 BUF_X1 output159 (.A(net170),
    .Z(data_addr_o[24]));
 BUF_X1 output160 (.A(net171),
    .Z(data_addr_o[25]));
 BUF_X1 output161 (.A(net172),
    .Z(data_addr_o[26]));
 BUF_X1 output162 (.A(net173),
    .Z(data_addr_o[27]));
 BUF_X1 output163 (.A(net174),
    .Z(data_addr_o[28]));
 BUF_X1 output164 (.A(net175),
    .Z(data_addr_o[29]));
 BUF_X1 output165 (.A(net176),
    .Z(data_addr_o[2]));
 BUF_X1 output166 (.A(net177),
    .Z(data_addr_o[30]));
 BUF_X1 output167 (.A(net178),
    .Z(data_addr_o[31]));
 BUF_X1 output168 (.A(net179),
    .Z(data_addr_o[3]));
 BUF_X1 output169 (.A(net180),
    .Z(data_addr_o[4]));
 BUF_X1 output170 (.A(net181),
    .Z(data_addr_o[5]));
 BUF_X1 output171 (.A(net182),
    .Z(data_addr_o[6]));
 BUF_X1 output172 (.A(net183),
    .Z(data_addr_o[7]));
 BUF_X1 output173 (.A(net184),
    .Z(data_addr_o[8]));
 BUF_X1 output174 (.A(net185),
    .Z(data_addr_o[9]));
 BUF_X1 output175 (.A(net186),
    .Z(data_be_o[0]));
 BUF_X1 output176 (.A(net187),
    .Z(data_be_o[1]));
 BUF_X1 output177 (.A(net188),
    .Z(data_be_o[2]));
 BUF_X1 output178 (.A(net189),
    .Z(data_be_o[3]));
 BUF_X1 output179 (.A(net190),
    .Z(data_req_o));
 BUF_X1 output180 (.A(net191),
    .Z(data_wdata_o[0]));
 BUF_X1 output181 (.A(net192),
    .Z(data_wdata_o[10]));
 BUF_X1 output182 (.A(net193),
    .Z(data_wdata_o[11]));
 BUF_X1 output183 (.A(net194),
    .Z(data_wdata_o[12]));
 BUF_X1 output184 (.A(net195),
    .Z(data_wdata_o[13]));
 BUF_X1 output185 (.A(net196),
    .Z(data_wdata_o[14]));
 BUF_X1 output186 (.A(net197),
    .Z(data_wdata_o[15]));
 BUF_X1 output187 (.A(net198),
    .Z(data_wdata_o[16]));
 BUF_X1 output188 (.A(net199),
    .Z(data_wdata_o[17]));
 BUF_X1 output189 (.A(net200),
    .Z(data_wdata_o[18]));
 BUF_X1 output190 (.A(net201),
    .Z(data_wdata_o[19]));
 BUF_X1 output191 (.A(net202),
    .Z(data_wdata_o[1]));
 BUF_X1 output192 (.A(net203),
    .Z(data_wdata_o[20]));
 BUF_X1 output193 (.A(net204),
    .Z(data_wdata_o[21]));
 BUF_X1 output194 (.A(net205),
    .Z(data_wdata_o[22]));
 BUF_X1 output195 (.A(net206),
    .Z(data_wdata_o[23]));
 BUF_X1 output196 (.A(net207),
    .Z(data_wdata_o[24]));
 BUF_X1 output197 (.A(net208),
    .Z(data_wdata_o[25]));
 BUF_X1 output198 (.A(net209),
    .Z(data_wdata_o[26]));
 BUF_X1 output199 (.A(net210),
    .Z(data_wdata_o[27]));
 BUF_X1 output200 (.A(net211),
    .Z(data_wdata_o[28]));
 BUF_X1 output201 (.A(net212),
    .Z(data_wdata_o[29]));
 BUF_X1 output202 (.A(net213),
    .Z(data_wdata_o[2]));
 BUF_X1 output203 (.A(net214),
    .Z(data_wdata_o[30]));
 BUF_X1 output204 (.A(net215),
    .Z(data_wdata_o[31]));
 BUF_X1 output205 (.A(net216),
    .Z(data_wdata_o[3]));
 BUF_X1 output206 (.A(net217),
    .Z(data_wdata_o[4]));
 BUF_X1 output207 (.A(net218),
    .Z(data_wdata_o[5]));
 BUF_X1 output208 (.A(net219),
    .Z(data_wdata_o[6]));
 BUF_X1 output209 (.A(net220),
    .Z(data_wdata_o[7]));
 BUF_X1 output210 (.A(net221),
    .Z(data_wdata_o[8]));
 BUF_X1 output211 (.A(net222),
    .Z(data_wdata_o[9]));
 BUF_X1 output212 (.A(net223),
    .Z(data_we_o));
 BUF_X1 output213 (.A(net224),
    .Z(instr_addr_o[10]));
 BUF_X1 output214 (.A(net225),
    .Z(instr_addr_o[11]));
 BUF_X1 output215 (.A(net226),
    .Z(instr_addr_o[12]));
 BUF_X1 output216 (.A(net227),
    .Z(instr_addr_o[13]));
 BUF_X1 output217 (.A(net228),
    .Z(instr_addr_o[14]));
 BUF_X1 output218 (.A(net229),
    .Z(instr_addr_o[15]));
 BUF_X1 output219 (.A(net230),
    .Z(instr_addr_o[16]));
 BUF_X1 output220 (.A(net231),
    .Z(instr_addr_o[17]));
 BUF_X1 output221 (.A(net232),
    .Z(instr_addr_o[18]));
 BUF_X1 output222 (.A(net233),
    .Z(instr_addr_o[19]));
 BUF_X1 output223 (.A(net234),
    .Z(instr_addr_o[20]));
 BUF_X1 output224 (.A(net235),
    .Z(instr_addr_o[21]));
 BUF_X1 output225 (.A(net236),
    .Z(instr_addr_o[22]));
 BUF_X1 output226 (.A(net237),
    .Z(instr_addr_o[23]));
 BUF_X1 output227 (.A(net238),
    .Z(instr_addr_o[24]));
 BUF_X1 output228 (.A(net239),
    .Z(instr_addr_o[25]));
 BUF_X1 output229 (.A(net240),
    .Z(instr_addr_o[26]));
 BUF_X1 output230 (.A(net241),
    .Z(instr_addr_o[27]));
 BUF_X1 output231 (.A(net242),
    .Z(instr_addr_o[28]));
 BUF_X1 output232 (.A(net243),
    .Z(instr_addr_o[29]));
 BUF_X1 output233 (.A(net244),
    .Z(instr_addr_o[2]));
 BUF_X1 output234 (.A(net245),
    .Z(instr_addr_o[30]));
 BUF_X1 output235 (.A(net246),
    .Z(instr_addr_o[31]));
 BUF_X1 output236 (.A(net247),
    .Z(instr_addr_o[3]));
 BUF_X1 output237 (.A(net248),
    .Z(instr_addr_o[4]));
 BUF_X1 output238 (.A(net249),
    .Z(instr_addr_o[5]));
 BUF_X1 output239 (.A(net250),
    .Z(instr_addr_o[6]));
 BUF_X1 output240 (.A(net251),
    .Z(instr_addr_o[7]));
 BUF_X1 output241 (.A(net252),
    .Z(instr_addr_o[8]));
 BUF_X1 output242 (.A(net253),
    .Z(instr_addr_o[9]));
 BUF_X1 output243 (.A(net254),
    .Z(instr_req_o));
 BUF_X32 wire244 (.A(net261),
    .Z(net255));
 BUF_X32 max_length245 (.A(net259),
    .Z(net256));
 BUF_X32 max_length246 (.A(net260),
    .Z(net257));
 BUF_X32 max_length247 (.A(net260),
    .Z(net258));
 BUF_X32 max_length248 (.A(net260),
    .Z(net259));
 BUF_X32 wire249 (.A(net261),
    .Z(net260));
 BUF_X32 max_length250 (.A(net262),
    .Z(net261));
 BUF_X32 max_length251 (.A(net153),
    .Z(net262));
 BUF_X32 max_length252 (.A(net264),
    .Z(net263));
 BUF_X32 max_length253 (.A(net265),
    .Z(net264));
 BUF_X32 max_length254 (.A(net153),
    .Z(net265));
 LOGIC0_X1 _29849__255 (.Z(net266));
 LOGIC0_X1 _29850__256 (.Z(net267));
 LOGIC0_X1 _29851__257 (.Z(net268));
 LOGIC0_X1 _29852__258 (.Z(net269));
 LOGIC0_X1 _29883__259 (.Z(net270));
 LOGIC0_X1 _29884__260 (.Z(net271));
 CLKBUF_X3 clkbuf_0_clk_i (.A(clk_i),
    .Z(clknet_0_clk_i));
 CLKBUF_X3 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_1_0__leaf_clk_i));
 CLKBUF_X3 clkbuf_leaf_0_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_0_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_1_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_1_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_2_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_2_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_3_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_3_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_4_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_4_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_5_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_5_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_6_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_6_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_7_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_7_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_8_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_8_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_9_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_9_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_10_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_10_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_11_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_11_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_12_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_12_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_13_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_13_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_14_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_14_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_15_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_15_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_16_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_16_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_17_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_17_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_18_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_18_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_19_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_19_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_20_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_20_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_21_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_21_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_22_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_22_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_23_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_23_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_24_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_24_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_25_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_25_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_26_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_26_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_27_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_27_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_28_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_28_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_29_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_29_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_30_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_30_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_31_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_31_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_32_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_32_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_33_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_33_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_34_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_34_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_35_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_35_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_36_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_36_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_37_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_37_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_38_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_38_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_39_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_39_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_40_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_40_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_41_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_41_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_42_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_42_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_43_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_43_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_44_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_44_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_45_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_45_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_46_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_46_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_47_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_47_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_48_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_48_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_49_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_49_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_50_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_50_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_51_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_51_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_52_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_52_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_53_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_53_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_54_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_54_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_55_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_55_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_56_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_56_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_57_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_57_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_58_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_58_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_59_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_59_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_60_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_60_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_61_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_61_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_62_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_62_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_63_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_63_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_64_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_64_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_65_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_65_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_66_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_66_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_67_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_67_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_68_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_68_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_69_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_69_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_70_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_70_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_71_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_71_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_72_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_72_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_73_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_73_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_74_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_74_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_75_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_75_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_76_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_76_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_77_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_77_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_78_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_78_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_79_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_79_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_80_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_80_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_81_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_81_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_82_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_82_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_83_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_83_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_84_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_84_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_85_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_85_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_86_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_86_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_87_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_87_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_88_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_88_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_89_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_89_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_90_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_90_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_91_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_91_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_92_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_92_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_93_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_93_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_94_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_94_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_95_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_95_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_96_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_96_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_97_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_97_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_98_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_98_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_99_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_99_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_100_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_100_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_101_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_101_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_102_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_102_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_103_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_103_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_104_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_104_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_105_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_105_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_106_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_106_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_107_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_107_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_108_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_108_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_109_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_109_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_110_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_110_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_111_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_111_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_112_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_112_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_113_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_113_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_114_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_114_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_115_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_115_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_116_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_116_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_117_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_117_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_118_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_118_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_119_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_119_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_120_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_120_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_121_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_121_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_122_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_122_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_123_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_123_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_124_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_124_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_125_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_125_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_126_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_126_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_127_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_127_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_128_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_128_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_129_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_129_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_130_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_130_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_131_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_131_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_132_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_132_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_133_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_133_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_134_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_134_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_135_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_135_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_136_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_136_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_137_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_137_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_138_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_138_clk_i_regs));
 CLKBUF_X3 clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .Z(clknet_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_0_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_0_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_1_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_1_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_2_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_2_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_3_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_3_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_4_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_4_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_5_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_5_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_6_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_6_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_7_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_7_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_8_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_8_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_9_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_9_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_10_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_10_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_11_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_11_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_12_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_12_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_13_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_13_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_14_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_14_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_15_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_15_0_clk_i_regs));
 INV_X2 clkload0 (.A(clknet_4_1_0_clk_i_regs));
 INV_X4 clkload1 (.A(clknet_4_3_0_clk_i_regs));
 INV_X4 clkload2 (.A(clknet_4_4_0_clk_i_regs));
 INV_X8 clkload3 (.A(clknet_4_5_0_clk_i_regs));
 INV_X2 clkload4 (.A(clknet_4_6_0_clk_i_regs));
 INV_X2 clkload5 (.A(clknet_4_7_0_clk_i_regs));
 CLKBUF_X3 clkload6 (.A(clknet_4_8_0_clk_i_regs));
 INV_X2 clkload7 (.A(clknet_4_9_0_clk_i_regs));
 INV_X2 clkload8 (.A(clknet_4_11_0_clk_i_regs));
 INV_X2 clkload9 (.A(clknet_4_12_0_clk_i_regs));
 INV_X2 clkload10 (.A(clknet_4_14_0_clk_i_regs));
 INV_X2 clkload11 (.A(clknet_4_15_0_clk_i_regs));
 CLKBUF_X1 clkload12 (.A(clknet_leaf_1_clk_i_regs));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_2_clk_i_regs));
 INV_X1 clkload14 (.A(clknet_leaf_4_clk_i_regs));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_7_clk_i_regs));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_135_clk_i_regs));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_137_clk_i_regs));
 INV_X1 clkload18 (.A(clknet_leaf_138_clk_i_regs));
 INV_X2 clkload19 (.A(clknet_leaf_123_clk_i_regs));
 INV_X1 clkload20 (.A(clknet_leaf_124_clk_i_regs));
 INV_X1 clkload21 (.A(clknet_leaf_129_clk_i_regs));
 INV_X1 clkload22 (.A(clknet_leaf_130_clk_i_regs));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_131_clk_i_regs));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_132_clk_i_regs));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_133_clk_i_regs));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_134_clk_i_regs));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_9_clk_i_regs));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_10_clk_i_regs));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_12_clk_i_regs));
 INV_X1 clkload30 (.A(clknet_leaf_14_clk_i_regs));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_15_clk_i_regs));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_16_clk_i_regs));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_33_clk_i_regs));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_18_clk_i_regs));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_20_clk_i_regs));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_125_clk_i_regs));
 INV_X1 clkload37 (.A(clknet_leaf_126_clk_i_regs));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_127_clk_i_regs));
 INV_X2 clkload39 (.A(clknet_leaf_107_clk_i_regs));
 INV_X2 clkload40 (.A(clknet_leaf_113_clk_i_regs));
 CLKBUF_X1 clkload41 (.A(clknet_leaf_21_clk_i_regs));
 INV_X1 clkload42 (.A(clknet_leaf_100_clk_i_regs));
 INV_X1 clkload43 (.A(clknet_leaf_116_clk_i_regs));
 INV_X1 clkload44 (.A(clknet_leaf_117_clk_i_regs));
 INV_X1 clkload45 (.A(clknet_leaf_118_clk_i_regs));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_120_clk_i_regs));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_121_clk_i_regs));
 INV_X2 clkload48 (.A(clknet_leaf_102_clk_i_regs));
 INV_X1 clkload49 (.A(clknet_leaf_103_clk_i_regs));
 INV_X1 clkload50 (.A(clknet_leaf_104_clk_i_regs));
 INV_X2 clkload51 (.A(clknet_leaf_105_clk_i_regs));
 INV_X2 clkload52 (.A(clknet_leaf_106_clk_i_regs));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_114_clk_i_regs));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_115_clk_i_regs));
 INV_X2 clkload55 (.A(clknet_leaf_29_clk_i_regs));
 INV_X2 clkload56 (.A(clknet_leaf_31_clk_i_regs));
 INV_X2 clkload57 (.A(clknet_leaf_32_clk_i_regs));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_34_clk_i_regs));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_35_clk_i_regs));
 INV_X2 clkload60 (.A(clknet_leaf_36_clk_i_regs));
 INV_X1 clkload61 (.A(clknet_leaf_38_clk_i_regs));
 INV_X1 clkload62 (.A(clknet_leaf_39_clk_i_regs));
 INV_X1 clkload63 (.A(clknet_leaf_40_clk_i_regs));
 CLKBUF_X1 clkload64 (.A(clknet_leaf_25_clk_i_regs));
 INV_X1 clkload65 (.A(clknet_leaf_27_clk_i_regs));
 CLKBUF_X1 clkload66 (.A(clknet_leaf_64_clk_i_regs));
 CLKBUF_X1 clkload67 (.A(clknet_leaf_65_clk_i_regs));
 CLKBUF_X1 clkload68 (.A(clknet_leaf_41_clk_i_regs));
 INV_X1 clkload69 (.A(clknet_leaf_43_clk_i_regs));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_44_clk_i_regs));
 CLKBUF_X1 clkload71 (.A(clknet_leaf_45_clk_i_regs));
 CLKBUF_X1 clkload72 (.A(clknet_leaf_49_clk_i_regs));
 CLKBUF_X1 clkload73 (.A(clknet_leaf_50_clk_i_regs));
 INV_X1 clkload74 (.A(clknet_leaf_51_clk_i_regs));
 CLKBUF_X1 clkload75 (.A(clknet_leaf_52_clk_i_regs));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_55_clk_i_regs));
 CLKBUF_X1 clkload77 (.A(clknet_leaf_59_clk_i_regs));
 CLKBUF_X1 clkload78 (.A(clknet_leaf_61_clk_i_regs));
 CLKBUF_X1 clkload79 (.A(clknet_leaf_62_clk_i_regs));
 CLKBUF_X1 clkload80 (.A(clknet_leaf_63_clk_i_regs));
 CLKBUF_X1 clkload81 (.A(clknet_leaf_22_clk_i_regs));
 CLKBUF_X1 clkload82 (.A(clknet_leaf_68_clk_i_regs));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_70_clk_i_regs));
 INV_X1 clkload84 (.A(clknet_leaf_72_clk_i_regs));
 CLKBUF_X1 clkload85 (.A(clknet_leaf_99_clk_i_regs));
 INV_X1 clkload86 (.A(clknet_leaf_89_clk_i_regs));
 CLKBUF_X1 clkload87 (.A(clknet_leaf_90_clk_i_regs));
 CLKBUF_X1 clkload88 (.A(clknet_leaf_92_clk_i_regs));
 CLKBUF_X1 clkload89 (.A(clknet_leaf_93_clk_i_regs));
 CLKBUF_X1 clkload90 (.A(clknet_leaf_95_clk_i_regs));
 CLKBUF_X1 clkload91 (.A(clknet_leaf_98_clk_i_regs));
 CLKBUF_X1 clkload92 (.A(clknet_leaf_57_clk_i_regs));
 CLKBUF_X1 clkload93 (.A(clknet_leaf_58_clk_i_regs));
 CLKBUF_X1 clkload94 (.A(clknet_leaf_75_clk_i_regs));
 INV_X1 clkload95 (.A(clknet_leaf_76_clk_i_regs));
 INV_X2 clkload96 (.A(clknet_leaf_77_clk_i_regs));
 CLKBUF_X1 clkload97 (.A(clknet_leaf_78_clk_i_regs));
 CLKBUF_X1 clkload98 (.A(clknet_leaf_79_clk_i_regs));
 INV_X1 clkload99 (.A(clknet_leaf_80_clk_i_regs));
 CLKBUF_X1 clkload100 (.A(clknet_leaf_74_clk_i_regs));
 CLKBUF_X1 clkload101 (.A(clknet_leaf_84_clk_i_regs));
 CLKBUF_X1 clkload102 (.A(clknet_leaf_85_clk_i_regs));
 CLKBUF_X1 clkload103 (.A(clknet_leaf_87_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X3 clkload104 (.A(clknet_4_0_0_clk));
 INV_X2 clkload105 (.A(clknet_4_1_0_clk));
 INV_X4 clkload106 (.A(clknet_4_2_0_clk));
 INV_X4 clkload107 (.A(clknet_4_3_0_clk));
 INV_X2 clkload108 (.A(clknet_4_4_0_clk));
 INV_X8 clkload109 (.A(clknet_4_6_0_clk));
 INV_X4 clkload110 (.A(clknet_4_7_0_clk));
 INV_X8 clkload111 (.A(clknet_4_8_0_clk));
 INV_X8 clkload112 (.A(clknet_4_9_0_clk));
 INV_X8 clkload113 (.A(clknet_4_10_0_clk));
 INV_X8 clkload114 (.A(clknet_4_11_0_clk));
 INV_X4 clkload115 (.A(clknet_4_12_0_clk));
 INV_X4 clkload116 (.A(clknet_4_13_0_clk));
 INV_X8 clkload117 (.A(clknet_4_14_0_clk));
 INV_X8 clkload118 (.A(clknet_4_15_0_clk));
 INV_X1 clkload119 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload120 (.A(clknet_leaf_1_clk));
 INV_X2 clkload121 (.A(clknet_leaf_127_clk));
 CLKBUF_X1 clkload122 (.A(clknet_leaf_128_clk));
 CLKBUF_X1 clkload123 (.A(clknet_leaf_129_clk));
 CLKBUF_X1 clkload124 (.A(clknet_leaf_130_clk));
 CLKBUF_X1 clkload125 (.A(clknet_leaf_133_clk));
 CLKBUF_X1 clkload126 (.A(clknet_leaf_135_clk));
 CLKBUF_X1 clkload127 (.A(clknet_leaf_102_clk));
 INV_X1 clkload128 (.A(clknet_leaf_104_clk));
 INV_X2 clkload129 (.A(clknet_leaf_118_clk));
 CLKBUF_X1 clkload130 (.A(clknet_leaf_119_clk));
 CLKBUF_X1 clkload131 (.A(clknet_leaf_120_clk));
 CLKBUF_X1 clkload132 (.A(clknet_leaf_121_clk));
 CLKBUF_X1 clkload133 (.A(clknet_leaf_123_clk));
 CLKBUF_X2 clkload134 (.A(clknet_leaf_125_clk));
 INV_X1 clkload135 (.A(clknet_leaf_126_clk));
 INV_X2 clkload136 (.A(clknet_leaf_2_clk));
 INV_X1 clkload137 (.A(clknet_leaf_3_clk));
 INV_X1 clkload138 (.A(clknet_leaf_4_clk));
 CLKBUF_X1 clkload139 (.A(clknet_leaf_5_clk));
 INV_X1 clkload140 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload141 (.A(clknet_leaf_7_clk));
 INV_X2 clkload142 (.A(clknet_leaf_9_clk));
 INV_X2 clkload143 (.A(clknet_leaf_109_clk));
 INV_X1 clkload144 (.A(clknet_leaf_110_clk));
 CLKBUF_X1 clkload145 (.A(clknet_leaf_111_clk));
 CLKBUF_X1 clkload146 (.A(clknet_leaf_112_clk));
 INV_X1 clkload147 (.A(clknet_leaf_113_clk));
 CLKBUF_X1 clkload148 (.A(clknet_leaf_115_clk));
 INV_X1 clkload149 (.A(clknet_leaf_117_clk));
 CLKBUF_X1 clkload150 (.A(clknet_leaf_94_clk));
 CLKBUF_X1 clkload151 (.A(clknet_leaf_96_clk));
 CLKBUF_X1 clkload152 (.A(clknet_leaf_97_clk));
 CLKBUF_X1 clkload153 (.A(clknet_leaf_98_clk));
 CLKBUF_X1 clkload154 (.A(clknet_leaf_99_clk));
 INV_X2 clkload155 (.A(clknet_leaf_100_clk));
 CLKBUF_X1 clkload156 (.A(clknet_leaf_101_clk));
 CLKBUF_X1 clkload157 (.A(clknet_leaf_103_clk));
 CLKBUF_X1 clkload158 (.A(clknet_leaf_105_clk));
 CLKBUF_X1 clkload159 (.A(clknet_leaf_106_clk));
 INV_X1 clkload160 (.A(clknet_leaf_80_clk));
 INV_X2 clkload161 (.A(clknet_leaf_81_clk));
 CLKBUF_X1 clkload162 (.A(clknet_leaf_82_clk));
 INV_X1 clkload163 (.A(clknet_leaf_83_clk));
 CLKBUF_X1 clkload164 (.A(clknet_leaf_84_clk));
 INV_X1 clkload165 (.A(clknet_leaf_85_clk));
 CLKBUF_X1 clkload166 (.A(clknet_leaf_86_clk));
 INV_X1 clkload167 (.A(clknet_leaf_87_clk));
 INV_X1 clkload168 (.A(clknet_leaf_88_clk));
 INV_X2 clkload169 (.A(clknet_leaf_89_clk));
 CLKBUF_X1 clkload170 (.A(clknet_leaf_90_clk));
 INV_X2 clkload171 (.A(clknet_leaf_91_clk));
 CLKBUF_X1 clkload172 (.A(clknet_leaf_92_clk));
 CLKBUF_X1 clkload173 (.A(clknet_leaf_59_clk));
 INV_X1 clkload174 (.A(clknet_leaf_60_clk));
 CLKBUF_X1 clkload175 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload176 (.A(clknet_leaf_62_clk));
 INV_X1 clkload177 (.A(clknet_leaf_107_clk));
 CLKBUF_X1 clkload178 (.A(clknet_leaf_108_clk));
 CLKBUF_X1 clkload179 (.A(clknet_leaf_64_clk));
 INV_X1 clkload180 (.A(clknet_leaf_65_clk));
 CLKBUF_X1 clkload181 (.A(clknet_leaf_72_clk));
 CLKBUF_X1 clkload182 (.A(clknet_leaf_73_clk));
 CLKBUF_X1 clkload183 (.A(clknet_leaf_74_clk));
 CLKBUF_X1 clkload184 (.A(clknet_leaf_75_clk));
 INV_X1 clkload185 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload186 (.A(clknet_leaf_77_clk));
 CLKBUF_X1 clkload187 (.A(clknet_leaf_79_clk));
 INV_X1 clkload188 (.A(clknet_leaf_10_clk));
 INV_X1 clkload189 (.A(clknet_leaf_11_clk));
 INV_X1 clkload190 (.A(clknet_leaf_19_clk));
 INV_X4 clkload191 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload192 (.A(clknet_leaf_12_clk));
 INV_X1 clkload193 (.A(clknet_leaf_14_clk));
 INV_X1 clkload194 (.A(clknet_leaf_15_clk));
 INV_X2 clkload195 (.A(clknet_leaf_18_clk));
 INV_X1 clkload196 (.A(clknet_leaf_24_clk));
 CLKBUF_X1 clkload197 (.A(clknet_leaf_26_clk));
 CLKBUF_X1 clkload198 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload199 (.A(clknet_leaf_31_clk));
 INV_X1 clkload200 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload201 (.A(clknet_leaf_23_clk));
 CLKBUF_X1 clkload202 (.A(clknet_leaf_28_clk));
 INV_X1 clkload203 (.A(clknet_leaf_53_clk));
 CLKBUF_X2 clkload204 (.A(clknet_leaf_49_clk));
 CLKBUF_X2 clkload205 (.A(clknet_leaf_50_clk));
 CLKBUF_X2 clkload206 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload207 (.A(clknet_leaf_54_clk));
 CLKBUF_X1 clkload208 (.A(clknet_leaf_55_clk));
 INV_X2 clkload209 (.A(clknet_leaf_57_clk));
 INV_X1 clkload210 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload211 (.A(clknet_leaf_66_clk));
 CLKBUF_X1 clkload212 (.A(clknet_leaf_44_clk));
 CLKBUF_X1 clkload213 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload214 (.A(clknet_leaf_46_clk));
 INV_X1 clkload215 (.A(clknet_leaf_47_clk));
 INV_X1 clkload216 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload217 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload218 (.A(clknet_leaf_69_clk));
 INV_X1 clkload219 (.A(clknet_leaf_70_clk));
 CLKBUF_X1 clkload220 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload221 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload222 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload223 (.A(clknet_leaf_34_clk));
 CLKBUF_X2 clkload224 (.A(clknet_leaf_35_clk));
 CLKBUF_X1 clkload225 (.A(clknet_leaf_36_clk));
 CLKBUF_X2 clkload226 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload227 (.A(clknet_leaf_38_clk));
 CLKBUF_X1 clkload228 (.A(clknet_leaf_39_clk));
 CLKBUF_X1 clkload229 (.A(clknet_leaf_40_clk));
 CLKBUF_X1 clkload230 (.A(clknet_leaf_41_clk));
 CLKBUF_X1 clkload231 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload232 (.A(clknet_leaf_43_clk));
 CLKBUF_X3 delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .Z(delaynet_1_core_clock));
 CLKBUF_X3 delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .Z(clk_i_regs));
 BUF_X1 rebuffer1 (.A(_03392_),
    .Z(net272));
 BUF_X1 rebuffer2 (.A(net272),
    .Z(net273));
 BUF_X1 rebuffer3 (.A(net272),
    .Z(net274));
 BUF_X1 rebuffer4 (.A(_03417_),
    .Z(net275));
 BUF_X1 rebuffer5 (.A(net275),
    .Z(net276));
 BUF_X2 rebuffer6 (.A(_10548_),
    .Z(net277));
 INV_X2 clone8 (.A(_03417_),
    .ZN(net279));
 BUF_X1 rebuffer9 (.A(net349),
    .Z(net280));
 BUF_X4 rebuffer10 (.A(net280),
    .Z(net281));
 BUF_X1 rebuffer11 (.A(_10511_),
    .Z(net282));
 BUF_X1 rebuffer12 (.A(net282),
    .Z(net283));
 BUF_X1 rebuffer13 (.A(net282),
    .Z(net284));
 BUF_X1 rebuffer14 (.A(net421),
    .Z(net285));
 BUF_X2 rebuffer15 (.A(net285),
    .Z(net286));
 BUF_X1 rebuffer16 (.A(_12823_),
    .Z(net287));
 BUF_X2 rebuffer17 (.A(net287),
    .Z(net288));
 BUF_X1 rebuffer18 (.A(_12725_),
    .Z(net289));
 BUF_X2 rebuffer19 (.A(net289),
    .Z(net290));
 MUX2_X1 clone20 (.A(_12144_),
    .B(_03275_),
    .S(_03655_),
    .Z(net291));
 BUF_X4 rebuffer22 (.A(_11470_),
    .Z(net293));
 BUF_X1 rebuffer23 (.A(net293),
    .Z(net294));
 BUF_X1 rebuffer24 (.A(net294),
    .Z(net295));
 BUF_X4 clone25 (.A(_12099_),
    .Z(net296));
 BUF_X1 rebuffer26 (.A(_15365_),
    .Z(net297));
 BUF_X1 rebuffer27 (.A(net297),
    .Z(net298));
 BUF_X8 clone29 (.A(_10310_),
    .Z(net300));
 BUF_X2 clone30 (.A(_15362_),
    .Z(net301));
 BUF_X1 rebuffer31 (.A(_10319_),
    .Z(net302));
 BUF_X1 rebuffer32 (.A(_11993_),
    .Z(net303));
 BUF_X8 clone33 (.A(_10310_),
    .Z(net304));
 BUF_X4 clone34 (.A(net306),
    .Z(net305));
 BUF_X1 rebuffer35 (.A(\id_stage_i.controller_i.instr_i[28] ),
    .Z(net306));
 BUF_X1 rebuffer36 (.A(_10332_),
    .Z(net307));
 BUF_X1 rebuffer37 (.A(net307),
    .Z(net308));
 BUF_X1 rebuffer38 (.A(net308),
    .Z(net309));
 BUF_X1 rebuffer39 (.A(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net310));
 BUF_X4 clone40 (.A(net312),
    .Z(net311));
 BUF_X1 rebuffer41 (.A(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net312));
 BUF_X2 rebuffer43 (.A(net313),
    .Z(net314));
 BUF_X4 clone44 (.A(net316),
    .Z(net315));
 BUF_X1 rebuffer45 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net316));
 BUF_X8 clone46 (.A(_04030_),
    .Z(net317));
 BUF_X2 rebuffer47 (.A(_15730_),
    .Z(net318));
 BUF_X4 rebuffer48 (.A(_11554_),
    .Z(net319));
 BUF_X1 rebuffer49 (.A(net319),
    .Z(net320));
 MUX2_X1 clone51 (.A(_11202_),
    .B(net421),
    .S(_03655_),
    .Z(net322));
 BUF_X4 clone52 (.A(_03703_),
    .Z(net323));
 MUX2_X1 clone53 (.A(_11158_),
    .B(_12823_),
    .S(_03655_),
    .Z(net324));
 BUF_X4 clone54 (.A(_03697_),
    .Z(net325));
 BUF_X32 clone55 (.A(_10459_),
    .Z(net326));
 BUF_X4 rebuffer56 (.A(_12221_),
    .Z(net327));
 BUF_X1 rebuffer57 (.A(_15700_),
    .Z(net328));
 BUF_X2 rebuffer58 (.A(_13224_),
    .Z(net329));
 BUF_X1 rebuffer59 (.A(_13314_),
    .Z(net330));
 BUF_X4 clone60 (.A(_04849_),
    .Z(net331));
 BUF_X4 clone61 (.A(_04849_),
    .Z(net332));
 BUF_X4 clone62 (.A(_04849_),
    .Z(net333));
 BUF_X8 clone63 (.A(_10335_),
    .Z(net334));
 BUF_X1 rebuffer64 (.A(net364),
    .Z(net335));
 BUF_X2 rebuffer65 (.A(_03717_),
    .Z(net336));
 BUF_X4 clone66 (.A(_03717_),
    .Z(net337));
 BUF_X4 clone67 (.A(_03676_),
    .Z(net338));
 MUX2_X1 clone68 (.A(_03675_),
    .B(_12392_),
    .S(_03656_),
    .Z(net339));
 BUF_X4 rebuffer69 (.A(_13258_),
    .Z(net340));
 BUF_X1 rebuffer70 (.A(net340),
    .Z(net341));
 BUF_X1 rebuffer71 (.A(net340),
    .Z(net342));
 BUF_X1 rebuffer72 (.A(net342),
    .Z(net343));
 AOI21_X2 clone73 (.A(_12374_),
    .B1(_10474_),
    .B2(_12391_),
    .ZN(net344));
 BUF_X1 rebuffer74 (.A(net348),
    .Z(net345));
 BUF_X4 rebuffer75 (.A(_12482_),
    .Z(net346));
 BUF_X4 rebuffer76 (.A(net346),
    .Z(net347));
 BUF_X4 rebuffer78 (.A(_12553_),
    .Z(net349));
 BUF_X4 rebuffer79 (.A(_13187_),
    .Z(net350));
 BUF_X1 rebuffer80 (.A(net350),
    .Z(net351));
 BUF_X1 rebuffer81 (.A(net350),
    .Z(net352));
 BUF_X1 rebuffer82 (.A(net352),
    .Z(net353));
 BUF_X4 clone83 (.A(_03661_),
    .Z(net354));
 BUF_X1 rebuffer84 (.A(_12651_),
    .Z(net355));
 BUF_X4 clone85 (.A(_05210_),
    .Z(net356));
 BUF_X16 clone86 (.A(_10457_),
    .Z(net357));
 BUF_X1 rebuffer89 (.A(net358),
    .Z(net360));
 BUF_X4 rebuffer90 (.A(_12757_),
    .Z(net361));
 BUF_X1 rebuffer91 (.A(net361),
    .Z(net362));
 BUF_X1 rebuffer92 (.A(net361),
    .Z(net363));
 BUF_X2 rebuffer94 (.A(_11398_),
    .Z(net365));
 XNOR2_X1 clone95 (.A(_12771_),
    .B(_12762_),
    .ZN(net366));
 BUF_X1 rebuffer96 (.A(net449),
    .Z(net367));
 BUF_X2 rebuffer97 (.A(net367),
    .Z(net368));
 BUF_X1 rebuffer98 (.A(\alu_adder_result_ex[18] ),
    .Z(net369));
 BUF_X1 rebuffer99 (.A(net369),
    .Z(net370));
 BUF_X1 rebuffer100 (.A(net370),
    .Z(net371));
 XNOR2_X1 clone101 (.A(_12944_),
    .B(_12937_),
    .ZN(net372));
 INV_X2 clone102 (.A(net374),
    .ZN(net373));
 BUF_X1 rebuffer103 (.A(_13111_),
    .Z(net374));
 BUF_X1 rebuffer104 (.A(\alu_adder_result_ex[27] ),
    .Z(net375));
 BUF_X1 rebuffer105 (.A(net375),
    .Z(net376));
 BUF_X1 rebuffer106 (.A(net375),
    .Z(net377));
 BUF_X4 rebuffer107 (.A(_08049_),
    .Z(net378));
 BUF_X2 rebuffer108 (.A(net378),
    .Z(net379));
 XNOR2_X1 clone109 (.A(_12280_),
    .B(_12262_),
    .ZN(net380));
 XNOR2_X1 clone110 (.A(_12600_),
    .B(_12592_),
    .ZN(net381));
 BUF_X1 rebuffer111 (.A(\alu_adder_result_ex[26] ),
    .Z(net382));
 BUF_X1 rebuffer112 (.A(net382),
    .Z(net383));
 BUF_X1 rebuffer113 (.A(net382),
    .Z(net384));
 BUF_X1 rebuffer114 (.A(net384),
    .Z(net385));
 XNOR2_X1 clone115 (.A(_11920_),
    .B(_11902_),
    .ZN(net386));
 CLKBUF_X1 hold116 (.A(rst_ni),
    .Z(net387));
 BUF_X4 clone26 (.A(_05210_),
    .Z(net392));
 BUF_X16 clone27 (.A(_10457_),
    .Z(net393));
 BUF_X16 clone35 (.A(_10456_),
    .Z(net397));
 BUF_X4 clone38 (.A(_05210_),
    .Z(net400));
 BUF_X16 clone39 (.A(_10456_),
    .Z(net401));
 BUF_X16 clone41 (.A(net430),
    .Z(net402));
 BUF_X2 clone42 (.A(_05973_),
    .Z(net403));
 BUF_X4 clone43 (.A(_06173_),
    .Z(net404));
 BUF_X4 clone45 (.A(_06173_),
    .Z(net405));
 BUF_X4 clone47 (.A(_06173_),
    .Z(net406));
 BUF_X4 clone56 (.A(_05093_),
    .Z(net408));
 BUF_X4 clone57 (.A(_05093_),
    .Z(net409));
 BUF_X4 clone58 (.A(_05093_),
    .Z(net410));
 BUF_X4 rebuffer60 (.A(_10813_),
    .Z(net411));
 BUF_X4 clone64 (.A(_04907_),
    .Z(net412));
 BUF_X1 rebuffer66 (.A(\alu_adder_result_ex[23] ),
    .Z(net413));
 BUF_X4 clone76 (.A(_05036_),
    .Z(net418));
 BUF_X4 clone78 (.A(_05036_),
    .Z(net419));
 BUF_X4 clone79 (.A(_04907_),
    .Z(net420));
 BUF_X4 rebuffer83 (.A(_12896_),
    .Z(net421));
 BUF_X8 clone84 (.A(_05259_),
    .Z(net422));
 BUF_X16 clone94 (.A(net430),
    .Z(net427));
 BUF_X16 clone96 (.A(net430),
    .Z(net428));
 BUF_X16 clone97 (.A(_11937_),
    .Z(net429));
 BUF_X32 clone98 (.A(_10459_),
    .Z(net430));
 MUX2_X1 clone99 (.A(_11898_),
    .B(net350),
    .S(_03664_),
    .Z(net431));
 BUF_X16 rebuffer101 (.A(_10335_),
    .Z(net432));
 BUF_X16 clone103 (.A(net437),
    .Z(net433));
 BUF_X16 clone104 (.A(net437),
    .Z(net434));
 BUF_X32 clone105 (.A(net326),
    .Z(net435));
 BUF_X16 clone106 (.A(net437),
    .Z(net436));
 BUF_X16 clone107 (.A(_10459_),
    .Z(net437));
 BUF_X8 clone108 (.A(_05259_),
    .Z(net438));
 BUF_X4 clone112 (.A(_05036_),
    .Z(net440));
 BUF_X8 clone113 (.A(_05259_),
    .Z(net441));
 BUF_X8 clone114 (.A(_04977_),
    .Z(net442));
 BUF_X16 clone117 (.A(_05147_),
    .Z(net444));
 BUF_X16 clone118 (.A(_05147_),
    .Z(net445));
 BUF_X16 clone120 (.A(_05147_),
    .Z(net447));
 BUF_X1 rebuffer121 (.A(_12432_),
    .Z(net448));
 BUF_X2 rebuffer122 (.A(_15418_),
    .Z(net449));
 BUF_X1 rebuffer123 (.A(\alu_adder_result_ex[18] ),
    .Z(net450));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X16 FILLER_0_385 ();
 FILLCELL_X8 FILLER_0_401 ();
 FILLCELL_X4 FILLER_0_409 ();
 FILLCELL_X2 FILLER_0_413 ();
 FILLCELL_X8 FILLER_0_439 ();
 FILLCELL_X4 FILLER_0_447 ();
 FILLCELL_X16 FILLER_0_458 ();
 FILLCELL_X2 FILLER_0_474 ();
 FILLCELL_X4 FILLER_0_482 ();
 FILLCELL_X2 FILLER_0_486 ();
 FILLCELL_X1 FILLER_0_488 ();
 FILLCELL_X2 FILLER_0_519 ();
 FILLCELL_X1 FILLER_0_521 ();
 FILLCELL_X1 FILLER_0_536 ();
 FILLCELL_X1 FILLER_0_545 ();
 FILLCELL_X1 FILLER_0_586 ();
 FILLCELL_X1 FILLER_0_605 ();
 FILLCELL_X1 FILLER_0_623 ();
 FILLCELL_X1 FILLER_0_645 ();
 FILLCELL_X2 FILLER_0_675 ();
 FILLCELL_X2 FILLER_0_680 ();
 FILLCELL_X1 FILLER_0_682 ();
 FILLCELL_X2 FILLER_0_689 ();
 FILLCELL_X4 FILLER_0_694 ();
 FILLCELL_X4 FILLER_0_701 ();
 FILLCELL_X4 FILLER_0_708 ();
 FILLCELL_X8 FILLER_0_715 ();
 FILLCELL_X2 FILLER_0_723 ();
 FILLCELL_X4 FILLER_0_747 ();
 FILLCELL_X2 FILLER_0_773 ();
 FILLCELL_X1 FILLER_0_775 ();
 FILLCELL_X1 FILLER_0_799 ();
 FILLCELL_X4 FILLER_0_824 ();
 FILLCELL_X2 FILLER_0_828 ();
 FILLCELL_X4 FILLER_0_834 ();
 FILLCELL_X2 FILLER_0_838 ();
 FILLCELL_X1 FILLER_0_843 ();
 FILLCELL_X1 FILLER_0_867 ();
 FILLCELL_X1 FILLER_0_872 ();
 FILLCELL_X8 FILLER_0_898 ();
 FILLCELL_X1 FILLER_0_906 ();
 FILLCELL_X16 FILLER_0_920 ();
 FILLCELL_X8 FILLER_0_956 ();
 FILLCELL_X4 FILLER_0_964 ();
 FILLCELL_X1 FILLER_0_968 ();
 FILLCELL_X1 FILLER_0_973 ();
 FILLCELL_X4 FILLER_0_994 ();
 FILLCELL_X2 FILLER_0_998 ();
 FILLCELL_X16 FILLER_0_1022 ();
 FILLCELL_X8 FILLER_0_1038 ();
 FILLCELL_X32 FILLER_0_1066 ();
 FILLCELL_X32 FILLER_0_1098 ();
 FILLCELL_X32 FILLER_0_1130 ();
 FILLCELL_X32 FILLER_0_1162 ();
 FILLCELL_X32 FILLER_0_1194 ();
 FILLCELL_X8 FILLER_0_1226 ();
 FILLCELL_X4 FILLER_0_1234 ();
 FILLCELL_X8 FILLER_0_1241 ();
 FILLCELL_X4 FILLER_0_1249 ();
 FILLCELL_X2 FILLER_0_1253 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X8 FILLER_1_417 ();
 FILLCELL_X4 FILLER_1_425 ();
 FILLCELL_X2 FILLER_1_429 ();
 FILLCELL_X1 FILLER_1_431 ();
 FILLCELL_X1 FILLER_1_456 ();
 FILLCELL_X1 FILLER_1_464 ();
 FILLCELL_X8 FILLER_1_482 ();
 FILLCELL_X2 FILLER_1_490 ();
 FILLCELL_X1 FILLER_1_492 ();
 FILLCELL_X1 FILLER_1_500 ();
 FILLCELL_X1 FILLER_1_508 ();
 FILLCELL_X1 FILLER_1_530 ();
 FILLCELL_X2 FILLER_1_548 ();
 FILLCELL_X2 FILLER_1_568 ();
 FILLCELL_X1 FILLER_1_610 ();
 FILLCELL_X1 FILLER_1_628 ();
 FILLCELL_X1 FILLER_1_632 ();
 FILLCELL_X1 FILLER_1_650 ();
 FILLCELL_X32 FILLER_1_658 ();
 FILLCELL_X16 FILLER_1_690 ();
 FILLCELL_X2 FILLER_1_706 ();
 FILLCELL_X8 FILLER_1_732 ();
 FILLCELL_X4 FILLER_1_740 ();
 FILLCELL_X1 FILLER_1_744 ();
 FILLCELL_X4 FILLER_1_749 ();
 FILLCELL_X1 FILLER_1_764 ();
 FILLCELL_X8 FILLER_1_771 ();
 FILLCELL_X1 FILLER_1_779 ();
 FILLCELL_X1 FILLER_1_788 ();
 FILLCELL_X2 FILLER_1_793 ();
 FILLCELL_X8 FILLER_1_800 ();
 FILLCELL_X2 FILLER_1_859 ();
 FILLCELL_X2 FILLER_1_864 ();
 FILLCELL_X1 FILLER_1_866 ();
 FILLCELL_X8 FILLER_1_911 ();
 FILLCELL_X4 FILLER_1_919 ();
 FILLCELL_X1 FILLER_1_923 ();
 FILLCELL_X4 FILLER_1_944 ();
 FILLCELL_X8 FILLER_1_1001 ();
 FILLCELL_X4 FILLER_1_1009 ();
 FILLCELL_X16 FILLER_1_1037 ();
 FILLCELL_X2 FILLER_1_1053 ();
 FILLCELL_X2 FILLER_1_1079 ();
 FILLCELL_X32 FILLER_1_1103 ();
 FILLCELL_X32 FILLER_1_1135 ();
 FILLCELL_X32 FILLER_1_1167 ();
 FILLCELL_X4 FILLER_1_1199 ();
 FILLCELL_X2 FILLER_1_1203 ();
 FILLCELL_X1 FILLER_1_1205 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X16 FILLER_2_385 ();
 FILLCELL_X8 FILLER_2_401 ();
 FILLCELL_X4 FILLER_2_409 ();
 FILLCELL_X2 FILLER_2_413 ();
 FILLCELL_X2 FILLER_2_453 ();
 FILLCELL_X4 FILLER_2_462 ();
 FILLCELL_X8 FILLER_2_473 ();
 FILLCELL_X4 FILLER_2_481 ();
 FILLCELL_X1 FILLER_2_485 ();
 FILLCELL_X4 FILLER_2_510 ();
 FILLCELL_X1 FILLER_2_514 ();
 FILLCELL_X4 FILLER_2_518 ();
 FILLCELL_X2 FILLER_2_522 ();
 FILLCELL_X2 FILLER_2_548 ();
 FILLCELL_X8 FILLER_2_580 ();
 FILLCELL_X2 FILLER_2_602 ();
 FILLCELL_X1 FILLER_2_604 ();
 FILLCELL_X2 FILLER_2_612 ();
 FILLCELL_X1 FILLER_2_614 ();
 FILLCELL_X1 FILLER_2_622 ();
 FILLCELL_X1 FILLER_2_630 ();
 FILLCELL_X8 FILLER_2_632 ();
 FILLCELL_X1 FILLER_2_640 ();
 FILLCELL_X32 FILLER_2_662 ();
 FILLCELL_X2 FILLER_2_719 ();
 FILLCELL_X4 FILLER_2_724 ();
 FILLCELL_X1 FILLER_2_731 ();
 FILLCELL_X2 FILLER_2_735 ();
 FILLCELL_X1 FILLER_2_750 ();
 FILLCELL_X2 FILLER_2_754 ();
 FILLCELL_X2 FILLER_2_760 ();
 FILLCELL_X2 FILLER_2_766 ();
 FILLCELL_X1 FILLER_2_768 ();
 FILLCELL_X8 FILLER_2_817 ();
 FILLCELL_X2 FILLER_2_825 ();
 FILLCELL_X8 FILLER_2_835 ();
 FILLCELL_X4 FILLER_2_843 ();
 FILLCELL_X2 FILLER_2_847 ();
 FILLCELL_X1 FILLER_2_849 ();
 FILLCELL_X8 FILLER_2_880 ();
 FILLCELL_X4 FILLER_2_888 ();
 FILLCELL_X2 FILLER_2_892 ();
 FILLCELL_X4 FILLER_2_903 ();
 FILLCELL_X1 FILLER_2_907 ();
 FILLCELL_X16 FILLER_2_924 ();
 FILLCELL_X4 FILLER_2_940 ();
 FILLCELL_X2 FILLER_2_944 ();
 FILLCELL_X1 FILLER_2_946 ();
 FILLCELL_X2 FILLER_2_963 ();
 FILLCELL_X4 FILLER_2_967 ();
 FILLCELL_X2 FILLER_2_971 ();
 FILLCELL_X1 FILLER_2_985 ();
 FILLCELL_X4 FILLER_2_1007 ();
 FILLCELL_X4 FILLER_2_1013 ();
 FILLCELL_X1 FILLER_2_1017 ();
 FILLCELL_X2 FILLER_2_1031 ();
 FILLCELL_X1 FILLER_2_1035 ();
 FILLCELL_X1 FILLER_2_1058 ();
 FILLCELL_X4 FILLER_2_1072 ();
 FILLCELL_X32 FILLER_2_1086 ();
 FILLCELL_X32 FILLER_2_1118 ();
 FILLCELL_X32 FILLER_2_1150 ();
 FILLCELL_X32 FILLER_2_1182 ();
 FILLCELL_X32 FILLER_2_1214 ();
 FILLCELL_X8 FILLER_2_1246 ();
 FILLCELL_X1 FILLER_2_1254 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X8 FILLER_3_417 ();
 FILLCELL_X2 FILLER_3_425 ();
 FILLCELL_X2 FILLER_3_434 ();
 FILLCELL_X1 FILLER_3_436 ();
 FILLCELL_X2 FILLER_3_454 ();
 FILLCELL_X4 FILLER_3_487 ();
 FILLCELL_X4 FILLER_3_525 ();
 FILLCELL_X2 FILLER_3_529 ();
 FILLCELL_X4 FILLER_3_548 ();
 FILLCELL_X2 FILLER_3_566 ();
 FILLCELL_X1 FILLER_3_568 ();
 FILLCELL_X2 FILLER_3_572 ();
 FILLCELL_X1 FILLER_3_574 ();
 FILLCELL_X2 FILLER_3_578 ();
 FILLCELL_X4 FILLER_3_641 ();
 FILLCELL_X2 FILLER_3_645 ();
 FILLCELL_X1 FILLER_3_647 ();
 FILLCELL_X32 FILLER_3_665 ();
 FILLCELL_X16 FILLER_3_697 ();
 FILLCELL_X4 FILLER_3_716 ();
 FILLCELL_X1 FILLER_3_727 ();
 FILLCELL_X1 FILLER_3_736 ();
 FILLCELL_X2 FILLER_3_741 ();
 FILLCELL_X1 FILLER_3_745 ();
 FILLCELL_X4 FILLER_3_760 ();
 FILLCELL_X2 FILLER_3_764 ();
 FILLCELL_X1 FILLER_3_766 ();
 FILLCELL_X4 FILLER_3_772 ();
 FILLCELL_X1 FILLER_3_776 ();
 FILLCELL_X4 FILLER_3_796 ();
 FILLCELL_X4 FILLER_3_809 ();
 FILLCELL_X2 FILLER_3_813 ();
 FILLCELL_X1 FILLER_3_815 ();
 FILLCELL_X8 FILLER_3_839 ();
 FILLCELL_X1 FILLER_3_857 ();
 FILLCELL_X1 FILLER_3_868 ();
 FILLCELL_X4 FILLER_3_906 ();
 FILLCELL_X2 FILLER_3_936 ();
 FILLCELL_X1 FILLER_3_938 ();
 FILLCELL_X4 FILLER_3_950 ();
 FILLCELL_X1 FILLER_3_954 ();
 FILLCELL_X1 FILLER_3_961 ();
 FILLCELL_X4 FILLER_3_983 ();
 FILLCELL_X1 FILLER_3_987 ();
 FILLCELL_X4 FILLER_3_990 ();
 FILLCELL_X2 FILLER_3_994 ();
 FILLCELL_X1 FILLER_3_996 ();
 FILLCELL_X1 FILLER_3_1004 ();
 FILLCELL_X4 FILLER_3_1016 ();
 FILLCELL_X1 FILLER_3_1050 ();
 FILLCELL_X1 FILLER_3_1063 ();
 FILLCELL_X1 FILLER_3_1070 ();
 FILLCELL_X32 FILLER_3_1115 ();
 FILLCELL_X32 FILLER_3_1147 ();
 FILLCELL_X32 FILLER_3_1179 ();
 FILLCELL_X32 FILLER_3_1211 ();
 FILLCELL_X8 FILLER_3_1243 ();
 FILLCELL_X4 FILLER_3_1251 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X16 FILLER_4_385 ();
 FILLCELL_X8 FILLER_4_401 ();
 FILLCELL_X4 FILLER_4_409 ();
 FILLCELL_X1 FILLER_4_413 ();
 FILLCELL_X8 FILLER_4_438 ();
 FILLCELL_X2 FILLER_4_475 ();
 FILLCELL_X2 FILLER_4_501 ();
 FILLCELL_X1 FILLER_4_510 ();
 FILLCELL_X4 FILLER_4_563 ();
 FILLCELL_X1 FILLER_4_589 ();
 FILLCELL_X8 FILLER_4_595 ();
 FILLCELL_X4 FILLER_4_603 ();
 FILLCELL_X1 FILLER_4_607 ();
 FILLCELL_X8 FILLER_4_620 ();
 FILLCELL_X2 FILLER_4_628 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X4 FILLER_4_632 ();
 FILLCELL_X2 FILLER_4_636 ();
 FILLCELL_X4 FILLER_4_645 ();
 FILLCELL_X8 FILLER_4_681 ();
 FILLCELL_X2 FILLER_4_689 ();
 FILLCELL_X1 FILLER_4_691 ();
 FILLCELL_X4 FILLER_4_712 ();
 FILLCELL_X1 FILLER_4_716 ();
 FILLCELL_X1 FILLER_4_721 ();
 FILLCELL_X1 FILLER_4_727 ();
 FILLCELL_X1 FILLER_4_732 ();
 FILLCELL_X2 FILLER_4_737 ();
 FILLCELL_X1 FILLER_4_739 ();
 FILLCELL_X2 FILLER_4_753 ();
 FILLCELL_X1 FILLER_4_755 ();
 FILLCELL_X4 FILLER_4_759 ();
 FILLCELL_X2 FILLER_4_763 ();
 FILLCELL_X1 FILLER_4_765 ();
 FILLCELL_X1 FILLER_4_776 ();
 FILLCELL_X4 FILLER_4_781 ();
 FILLCELL_X1 FILLER_4_785 ();
 FILLCELL_X1 FILLER_4_798 ();
 FILLCELL_X2 FILLER_4_810 ();
 FILLCELL_X4 FILLER_4_835 ();
 FILLCELL_X1 FILLER_4_848 ();
 FILLCELL_X1 FILLER_4_857 ();
 FILLCELL_X1 FILLER_4_862 ();
 FILLCELL_X2 FILLER_4_871 ();
 FILLCELL_X1 FILLER_4_873 ();
 FILLCELL_X16 FILLER_4_882 ();
 FILLCELL_X2 FILLER_4_898 ();
 FILLCELL_X2 FILLER_4_909 ();
 FILLCELL_X1 FILLER_4_911 ();
 FILLCELL_X4 FILLER_4_921 ();
 FILLCELL_X2 FILLER_4_925 ();
 FILLCELL_X1 FILLER_4_961 ();
 FILLCELL_X2 FILLER_4_975 ();
 FILLCELL_X1 FILLER_4_977 ();
 FILLCELL_X1 FILLER_4_985 ();
 FILLCELL_X1 FILLER_4_994 ();
 FILLCELL_X2 FILLER_4_1002 ();
 FILLCELL_X4 FILLER_4_1026 ();
 FILLCELL_X1 FILLER_4_1030 ();
 FILLCELL_X2 FILLER_4_1036 ();
 FILLCELL_X1 FILLER_4_1046 ();
 FILLCELL_X1 FILLER_4_1049 ();
 FILLCELL_X1 FILLER_4_1054 ();
 FILLCELL_X8 FILLER_4_1062 ();
 FILLCELL_X4 FILLER_4_1070 ();
 FILLCELL_X2 FILLER_4_1074 ();
 FILLCELL_X32 FILLER_4_1095 ();
 FILLCELL_X32 FILLER_4_1127 ();
 FILLCELL_X32 FILLER_4_1159 ();
 FILLCELL_X32 FILLER_4_1191 ();
 FILLCELL_X32 FILLER_4_1223 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X16 FILLER_5_385 ();
 FILLCELL_X1 FILLER_5_401 ();
 FILLCELL_X8 FILLER_5_419 ();
 FILLCELL_X4 FILLER_5_427 ();
 FILLCELL_X2 FILLER_5_431 ();
 FILLCELL_X16 FILLER_5_445 ();
 FILLCELL_X2 FILLER_5_461 ();
 FILLCELL_X16 FILLER_5_470 ();
 FILLCELL_X2 FILLER_5_486 ();
 FILLCELL_X1 FILLER_5_495 ();
 FILLCELL_X4 FILLER_5_520 ();
 FILLCELL_X2 FILLER_5_534 ();
 FILLCELL_X1 FILLER_5_536 ();
 FILLCELL_X8 FILLER_5_542 ();
 FILLCELL_X1 FILLER_5_550 ();
 FILLCELL_X8 FILLER_5_558 ();
 FILLCELL_X2 FILLER_5_566 ();
 FILLCELL_X4 FILLER_5_582 ();
 FILLCELL_X1 FILLER_5_586 ();
 FILLCELL_X2 FILLER_5_604 ();
 FILLCELL_X16 FILLER_5_623 ();
 FILLCELL_X8 FILLER_5_639 ();
 FILLCELL_X4 FILLER_5_647 ();
 FILLCELL_X2 FILLER_5_651 ();
 FILLCELL_X1 FILLER_5_653 ();
 FILLCELL_X8 FILLER_5_678 ();
 FILLCELL_X4 FILLER_5_686 ();
 FILLCELL_X1 FILLER_5_690 ();
 FILLCELL_X8 FILLER_5_717 ();
 FILLCELL_X4 FILLER_5_725 ();
 FILLCELL_X2 FILLER_5_729 ();
 FILLCELL_X1 FILLER_5_731 ();
 FILLCELL_X1 FILLER_5_737 ();
 FILLCELL_X2 FILLER_5_745 ();
 FILLCELL_X1 FILLER_5_756 ();
 FILLCELL_X2 FILLER_5_775 ();
 FILLCELL_X8 FILLER_5_789 ();
 FILLCELL_X1 FILLER_5_797 ();
 FILLCELL_X1 FILLER_5_817 ();
 FILLCELL_X4 FILLER_5_836 ();
 FILLCELL_X2 FILLER_5_840 ();
 FILLCELL_X2 FILLER_5_851 ();
 FILLCELL_X8 FILLER_5_890 ();
 FILLCELL_X2 FILLER_5_898 ();
 FILLCELL_X16 FILLER_5_917 ();
 FILLCELL_X8 FILLER_5_933 ();
 FILLCELL_X8 FILLER_5_945 ();
 FILLCELL_X4 FILLER_5_953 ();
 FILLCELL_X1 FILLER_5_957 ();
 FILLCELL_X4 FILLER_5_960 ();
 FILLCELL_X8 FILLER_5_983 ();
 FILLCELL_X2 FILLER_5_991 ();
 FILLCELL_X1 FILLER_5_993 ();
 FILLCELL_X8 FILLER_5_1001 ();
 FILLCELL_X1 FILLER_5_1009 ();
 FILLCELL_X1 FILLER_5_1015 ();
 FILLCELL_X1 FILLER_5_1024 ();
 FILLCELL_X2 FILLER_5_1032 ();
 FILLCELL_X1 FILLER_5_1034 ();
 FILLCELL_X1 FILLER_5_1040 ();
 FILLCELL_X2 FILLER_5_1054 ();
 FILLCELL_X1 FILLER_5_1056 ();
 FILLCELL_X2 FILLER_5_1064 ();
 FILLCELL_X1 FILLER_5_1080 ();
 FILLCELL_X2 FILLER_5_1093 ();
 FILLCELL_X1 FILLER_5_1095 ();
 FILLCELL_X8 FILLER_5_1118 ();
 FILLCELL_X4 FILLER_5_1126 ();
 FILLCELL_X1 FILLER_5_1130 ();
 FILLCELL_X32 FILLER_5_1134 ();
 FILLCELL_X32 FILLER_5_1166 ();
 FILLCELL_X32 FILLER_5_1198 ();
 FILLCELL_X16 FILLER_5_1230 ();
 FILLCELL_X8 FILLER_5_1246 ();
 FILLCELL_X1 FILLER_5_1254 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X16 FILLER_6_353 ();
 FILLCELL_X8 FILLER_6_369 ();
 FILLCELL_X4 FILLER_6_377 ();
 FILLCELL_X2 FILLER_6_398 ();
 FILLCELL_X1 FILLER_6_400 ();
 FILLCELL_X8 FILLER_6_408 ();
 FILLCELL_X4 FILLER_6_416 ();
 FILLCELL_X1 FILLER_6_451 ();
 FILLCELL_X4 FILLER_6_469 ();
 FILLCELL_X4 FILLER_6_497 ();
 FILLCELL_X2 FILLER_6_501 ();
 FILLCELL_X1 FILLER_6_503 ();
 FILLCELL_X1 FILLER_6_512 ();
 FILLCELL_X8 FILLER_6_537 ();
 FILLCELL_X2 FILLER_6_545 ();
 FILLCELL_X4 FILLER_6_571 ();
 FILLCELL_X4 FILLER_6_582 ();
 FILLCELL_X2 FILLER_6_586 ();
 FILLCELL_X4 FILLER_6_602 ();
 FILLCELL_X1 FILLER_6_613 ();
 FILLCELL_X2 FILLER_6_632 ();
 FILLCELL_X1 FILLER_6_646 ();
 FILLCELL_X1 FILLER_6_659 ();
 FILLCELL_X16 FILLER_6_667 ();
 FILLCELL_X1 FILLER_6_683 ();
 FILLCELL_X8 FILLER_6_709 ();
 FILLCELL_X2 FILLER_6_735 ();
 FILLCELL_X1 FILLER_6_737 ();
 FILLCELL_X16 FILLER_6_750 ();
 FILLCELL_X4 FILLER_6_766 ();
 FILLCELL_X1 FILLER_6_770 ();
 FILLCELL_X2 FILLER_6_778 ();
 FILLCELL_X4 FILLER_6_789 ();
 FILLCELL_X2 FILLER_6_798 ();
 FILLCELL_X8 FILLER_6_817 ();
 FILLCELL_X1 FILLER_6_825 ();
 FILLCELL_X8 FILLER_6_830 ();
 FILLCELL_X2 FILLER_6_873 ();
 FILLCELL_X8 FILLER_6_893 ();
 FILLCELL_X4 FILLER_6_901 ();
 FILLCELL_X2 FILLER_6_905 ();
 FILLCELL_X1 FILLER_6_907 ();
 FILLCELL_X2 FILLER_6_970 ();
 FILLCELL_X1 FILLER_6_972 ();
 FILLCELL_X1 FILLER_6_975 ();
 FILLCELL_X1 FILLER_6_979 ();
 FILLCELL_X1 FILLER_6_985 ();
 FILLCELL_X1 FILLER_6_990 ();
 FILLCELL_X1 FILLER_6_995 ();
 FILLCELL_X2 FILLER_6_1000 ();
 FILLCELL_X8 FILLER_6_1006 ();
 FILLCELL_X2 FILLER_6_1014 ();
 FILLCELL_X8 FILLER_6_1046 ();
 FILLCELL_X4 FILLER_6_1054 ();
 FILLCELL_X8 FILLER_6_1066 ();
 FILLCELL_X1 FILLER_6_1088 ();
 FILLCELL_X2 FILLER_6_1092 ();
 FILLCELL_X32 FILLER_6_1140 ();
 FILLCELL_X16 FILLER_6_1172 ();
 FILLCELL_X8 FILLER_6_1188 ();
 FILLCELL_X4 FILLER_6_1196 ();
 FILLCELL_X2 FILLER_6_1200 ();
 FILLCELL_X1 FILLER_6_1206 ();
 FILLCELL_X32 FILLER_6_1210 ();
 FILLCELL_X8 FILLER_6_1242 ();
 FILLCELL_X4 FILLER_6_1250 ();
 FILLCELL_X1 FILLER_6_1254 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X4 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_403 ();
 FILLCELL_X1 FILLER_7_405 ();
 FILLCELL_X16 FILLER_7_419 ();
 FILLCELL_X1 FILLER_7_442 ();
 FILLCELL_X1 FILLER_7_460 ();
 FILLCELL_X2 FILLER_7_468 ();
 FILLCELL_X4 FILLER_7_494 ();
 FILLCELL_X1 FILLER_7_498 ();
 FILLCELL_X1 FILLER_7_516 ();
 FILLCELL_X4 FILLER_7_524 ();
 FILLCELL_X16 FILLER_7_535 ();
 FILLCELL_X8 FILLER_7_558 ();
 FILLCELL_X2 FILLER_7_566 ();
 FILLCELL_X8 FILLER_7_585 ();
 FILLCELL_X2 FILLER_7_593 ();
 FILLCELL_X1 FILLER_7_595 ();
 FILLCELL_X2 FILLER_7_603 ();
 FILLCELL_X2 FILLER_7_629 ();
 FILLCELL_X4 FILLER_7_638 ();
 FILLCELL_X1 FILLER_7_642 ();
 FILLCELL_X1 FILLER_7_672 ();
 FILLCELL_X2 FILLER_7_698 ();
 FILLCELL_X2 FILLER_7_722 ();
 FILLCELL_X2 FILLER_7_736 ();
 FILLCELL_X1 FILLER_7_738 ();
 FILLCELL_X1 FILLER_7_756 ();
 FILLCELL_X4 FILLER_7_797 ();
 FILLCELL_X1 FILLER_7_801 ();
 FILLCELL_X2 FILLER_7_806 ();
 FILLCELL_X1 FILLER_7_808 ();
 FILLCELL_X16 FILLER_7_811 ();
 FILLCELL_X2 FILLER_7_827 ();
 FILLCELL_X2 FILLER_7_834 ();
 FILLCELL_X1 FILLER_7_836 ();
 FILLCELL_X8 FILLER_7_844 ();
 FILLCELL_X2 FILLER_7_852 ();
 FILLCELL_X4 FILLER_7_866 ();
 FILLCELL_X2 FILLER_7_870 ();
 FILLCELL_X8 FILLER_7_879 ();
 FILLCELL_X4 FILLER_7_887 ();
 FILLCELL_X2 FILLER_7_891 ();
 FILLCELL_X1 FILLER_7_893 ();
 FILLCELL_X2 FILLER_7_942 ();
 FILLCELL_X1 FILLER_7_944 ();
 FILLCELL_X4 FILLER_7_949 ();
 FILLCELL_X16 FILLER_7_963 ();
 FILLCELL_X8 FILLER_7_979 ();
 FILLCELL_X4 FILLER_7_987 ();
 FILLCELL_X2 FILLER_7_991 ();
 FILLCELL_X1 FILLER_7_993 ();
 FILLCELL_X4 FILLER_7_1018 ();
 FILLCELL_X2 FILLER_7_1022 ();
 FILLCELL_X1 FILLER_7_1024 ();
 FILLCELL_X16 FILLER_7_1032 ();
 FILLCELL_X2 FILLER_7_1048 ();
 FILLCELL_X2 FILLER_7_1060 ();
 FILLCELL_X1 FILLER_7_1062 ();
 FILLCELL_X2 FILLER_7_1066 ();
 FILLCELL_X2 FILLER_7_1077 ();
 FILLCELL_X1 FILLER_7_1079 ();
 FILLCELL_X2 FILLER_7_1083 ();
 FILLCELL_X16 FILLER_7_1128 ();
 FILLCELL_X8 FILLER_7_1144 ();
 FILLCELL_X4 FILLER_7_1152 ();
 FILLCELL_X2 FILLER_7_1156 ();
 FILLCELL_X1 FILLER_7_1158 ();
 FILLCELL_X4 FILLER_7_1163 ();
 FILLCELL_X8 FILLER_7_1170 ();
 FILLCELL_X4 FILLER_7_1178 ();
 FILLCELL_X1 FILLER_7_1182 ();
 FILLCELL_X2 FILLER_7_1187 ();
 FILLCELL_X1 FILLER_7_1189 ();
 FILLCELL_X4 FILLER_7_1193 ();
 FILLCELL_X1 FILLER_7_1197 ();
 FILLCELL_X32 FILLER_7_1218 ();
 FILLCELL_X4 FILLER_7_1250 ();
 FILLCELL_X1 FILLER_7_1254 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X16 FILLER_8_353 ();
 FILLCELL_X8 FILLER_8_369 ();
 FILLCELL_X4 FILLER_8_384 ();
 FILLCELL_X2 FILLER_8_410 ();
 FILLCELL_X4 FILLER_8_419 ();
 FILLCELL_X2 FILLER_8_423 ();
 FILLCELL_X1 FILLER_8_425 ();
 FILLCELL_X4 FILLER_8_433 ();
 FILLCELL_X1 FILLER_8_437 ();
 FILLCELL_X8 FILLER_8_452 ();
 FILLCELL_X4 FILLER_8_460 ();
 FILLCELL_X2 FILLER_8_464 ();
 FILLCELL_X1 FILLER_8_478 ();
 FILLCELL_X4 FILLER_8_486 ();
 FILLCELL_X8 FILLER_8_497 ();
 FILLCELL_X4 FILLER_8_505 ();
 FILLCELL_X2 FILLER_8_516 ();
 FILLCELL_X4 FILLER_8_542 ();
 FILLCELL_X4 FILLER_8_570 ();
 FILLCELL_X4 FILLER_8_581 ();
 FILLCELL_X1 FILLER_8_585 ();
 FILLCELL_X4 FILLER_8_603 ();
 FILLCELL_X1 FILLER_8_607 ();
 FILLCELL_X16 FILLER_8_615 ();
 FILLCELL_X2 FILLER_8_632 ();
 FILLCELL_X4 FILLER_8_658 ();
 FILLCELL_X16 FILLER_8_669 ();
 FILLCELL_X8 FILLER_8_685 ();
 FILLCELL_X1 FILLER_8_693 ();
 FILLCELL_X2 FILLER_8_698 ();
 FILLCELL_X1 FILLER_8_700 ();
 FILLCELL_X8 FILLER_8_706 ();
 FILLCELL_X4 FILLER_8_714 ();
 FILLCELL_X1 FILLER_8_718 ();
 FILLCELL_X2 FILLER_8_745 ();
 FILLCELL_X2 FILLER_8_751 ();
 FILLCELL_X4 FILLER_8_774 ();
 FILLCELL_X1 FILLER_8_778 ();
 FILLCELL_X16 FILLER_8_787 ();
 FILLCELL_X1 FILLER_8_803 ();
 FILLCELL_X2 FILLER_8_808 ();
 FILLCELL_X2 FILLER_8_821 ();
 FILLCELL_X1 FILLER_8_823 ();
 FILLCELL_X2 FILLER_8_844 ();
 FILLCELL_X1 FILLER_8_869 ();
 FILLCELL_X8 FILLER_8_890 ();
 FILLCELL_X4 FILLER_8_898 ();
 FILLCELL_X1 FILLER_8_902 ();
 FILLCELL_X8 FILLER_8_921 ();
 FILLCELL_X2 FILLER_8_929 ();
 FILLCELL_X1 FILLER_8_931 ();
 FILLCELL_X1 FILLER_8_939 ();
 FILLCELL_X2 FILLER_8_953 ();
 FILLCELL_X1 FILLER_8_959 ();
 FILLCELL_X1 FILLER_8_964 ();
 FILLCELL_X4 FILLER_8_996 ();
 FILLCELL_X2 FILLER_8_1000 ();
 FILLCELL_X2 FILLER_8_1023 ();
 FILLCELL_X2 FILLER_8_1039 ();
 FILLCELL_X8 FILLER_8_1094 ();
 FILLCELL_X2 FILLER_8_1102 ();
 FILLCELL_X1 FILLER_8_1104 ();
 FILLCELL_X4 FILLER_8_1112 ();
 FILLCELL_X2 FILLER_8_1116 ();
 FILLCELL_X4 FILLER_8_1145 ();
 FILLCELL_X1 FILLER_8_1149 ();
 FILLCELL_X1 FILLER_8_1170 ();
 FILLCELL_X2 FILLER_8_1175 ();
 FILLCELL_X2 FILLER_8_1180 ();
 FILLCELL_X32 FILLER_8_1205 ();
 FILLCELL_X16 FILLER_8_1237 ();
 FILLCELL_X2 FILLER_8_1253 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X8 FILLER_9_353 ();
 FILLCELL_X4 FILLER_9_361 ();
 FILLCELL_X2 FILLER_9_396 ();
 FILLCELL_X1 FILLER_9_398 ();
 FILLCELL_X8 FILLER_9_423 ();
 FILLCELL_X4 FILLER_9_431 ();
 FILLCELL_X2 FILLER_9_435 ();
 FILLCELL_X2 FILLER_9_461 ();
 FILLCELL_X1 FILLER_9_463 ();
 FILLCELL_X8 FILLER_9_502 ();
 FILLCELL_X2 FILLER_9_510 ();
 FILLCELL_X1 FILLER_9_512 ();
 FILLCELL_X8 FILLER_9_541 ();
 FILLCELL_X2 FILLER_9_556 ();
 FILLCELL_X2 FILLER_9_565 ();
 FILLCELL_X1 FILLER_9_567 ();
 FILLCELL_X2 FILLER_9_585 ();
 FILLCELL_X1 FILLER_9_587 ();
 FILLCELL_X4 FILLER_9_602 ();
 FILLCELL_X4 FILLER_9_613 ();
 FILLCELL_X2 FILLER_9_624 ();
 FILLCELL_X1 FILLER_9_626 ();
 FILLCELL_X4 FILLER_9_651 ();
 FILLCELL_X16 FILLER_9_662 ();
 FILLCELL_X1 FILLER_9_678 ();
 FILLCELL_X1 FILLER_9_699 ();
 FILLCELL_X2 FILLER_9_731 ();
 FILLCELL_X1 FILLER_9_733 ();
 FILLCELL_X2 FILLER_9_745 ();
 FILLCELL_X1 FILLER_9_747 ();
 FILLCELL_X1 FILLER_9_752 ();
 FILLCELL_X16 FILLER_9_765 ();
 FILLCELL_X8 FILLER_9_781 ();
 FILLCELL_X1 FILLER_9_789 ();
 FILLCELL_X4 FILLER_9_795 ();
 FILLCELL_X4 FILLER_9_804 ();
 FILLCELL_X1 FILLER_9_812 ();
 FILLCELL_X1 FILLER_9_817 ();
 FILLCELL_X4 FILLER_9_822 ();
 FILLCELL_X2 FILLER_9_826 ();
 FILLCELL_X1 FILLER_9_828 ();
 FILLCELL_X1 FILLER_9_864 ();
 FILLCELL_X2 FILLER_9_873 ();
 FILLCELL_X4 FILLER_9_895 ();
 FILLCELL_X2 FILLER_9_908 ();
 FILLCELL_X4 FILLER_9_919 ();
 FILLCELL_X1 FILLER_9_945 ();
 FILLCELL_X2 FILLER_9_950 ();
 FILLCELL_X1 FILLER_9_955 ();
 FILLCELL_X2 FILLER_9_960 ();
 FILLCELL_X1 FILLER_9_967 ();
 FILLCELL_X4 FILLER_9_972 ();
 FILLCELL_X2 FILLER_9_976 ();
 FILLCELL_X1 FILLER_9_978 ();
 FILLCELL_X1 FILLER_9_989 ();
 FILLCELL_X8 FILLER_9_995 ();
 FILLCELL_X4 FILLER_9_1003 ();
 FILLCELL_X2 FILLER_9_1007 ();
 FILLCELL_X1 FILLER_9_1009 ();
 FILLCELL_X2 FILLER_9_1054 ();
 FILLCELL_X16 FILLER_9_1064 ();
 FILLCELL_X8 FILLER_9_1080 ();
 FILLCELL_X4 FILLER_9_1088 ();
 FILLCELL_X2 FILLER_9_1092 ();
 FILLCELL_X4 FILLER_9_1100 ();
 FILLCELL_X2 FILLER_9_1104 ();
 FILLCELL_X1 FILLER_9_1106 ();
 FILLCELL_X8 FILLER_9_1110 ();
 FILLCELL_X1 FILLER_9_1118 ();
 FILLCELL_X2 FILLER_9_1199 ();
 FILLCELL_X16 FILLER_9_1225 ();
 FILLCELL_X8 FILLER_9_1241 ();
 FILLCELL_X4 FILLER_9_1249 ();
 FILLCELL_X2 FILLER_9_1253 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X8 FILLER_10_385 ();
 FILLCELL_X2 FILLER_10_393 ();
 FILLCELL_X1 FILLER_10_395 ();
 FILLCELL_X4 FILLER_10_420 ();
 FILLCELL_X2 FILLER_10_424 ();
 FILLCELL_X1 FILLER_10_426 ();
 FILLCELL_X2 FILLER_10_441 ();
 FILLCELL_X8 FILLER_10_457 ();
 FILLCELL_X4 FILLER_10_465 ();
 FILLCELL_X1 FILLER_10_469 ();
 FILLCELL_X8 FILLER_10_477 ();
 FILLCELL_X1 FILLER_10_485 ();
 FILLCELL_X2 FILLER_10_491 ();
 FILLCELL_X2 FILLER_10_496 ();
 FILLCELL_X1 FILLER_10_498 ();
 FILLCELL_X2 FILLER_10_506 ();
 FILLCELL_X4 FILLER_10_513 ();
 FILLCELL_X1 FILLER_10_530 ();
 FILLCELL_X1 FILLER_10_538 ();
 FILLCELL_X8 FILLER_10_563 ();
 FILLCELL_X1 FILLER_10_571 ();
 FILLCELL_X1 FILLER_10_579 ();
 FILLCELL_X1 FILLER_10_587 ();
 FILLCELL_X1 FILLER_10_595 ();
 FILLCELL_X2 FILLER_10_603 ();
 FILLCELL_X4 FILLER_10_626 ();
 FILLCELL_X1 FILLER_10_630 ();
 FILLCELL_X16 FILLER_10_632 ();
 FILLCELL_X1 FILLER_10_648 ();
 FILLCELL_X2 FILLER_10_663 ();
 FILLCELL_X1 FILLER_10_665 ();
 FILLCELL_X4 FILLER_10_686 ();
 FILLCELL_X2 FILLER_10_690 ();
 FILLCELL_X1 FILLER_10_692 ();
 FILLCELL_X4 FILLER_10_697 ();
 FILLCELL_X8 FILLER_10_706 ();
 FILLCELL_X4 FILLER_10_714 ();
 FILLCELL_X2 FILLER_10_718 ();
 FILLCELL_X2 FILLER_10_746 ();
 FILLCELL_X2 FILLER_10_760 ();
 FILLCELL_X1 FILLER_10_762 ();
 FILLCELL_X8 FILLER_10_767 ();
 FILLCELL_X4 FILLER_10_775 ();
 FILLCELL_X1 FILLER_10_779 ();
 FILLCELL_X2 FILLER_10_823 ();
 FILLCELL_X1 FILLER_10_825 ();
 FILLCELL_X2 FILLER_10_829 ();
 FILLCELL_X1 FILLER_10_831 ();
 FILLCELL_X2 FILLER_10_836 ();
 FILLCELL_X1 FILLER_10_838 ();
 FILLCELL_X2 FILLER_10_842 ();
 FILLCELL_X2 FILLER_10_850 ();
 FILLCELL_X2 FILLER_10_862 ();
 FILLCELL_X1 FILLER_10_864 ();
 FILLCELL_X2 FILLER_10_869 ();
 FILLCELL_X8 FILLER_10_880 ();
 FILLCELL_X2 FILLER_10_888 ();
 FILLCELL_X8 FILLER_10_897 ();
 FILLCELL_X2 FILLER_10_905 ();
 FILLCELL_X1 FILLER_10_907 ();
 FILLCELL_X8 FILLER_10_917 ();
 FILLCELL_X4 FILLER_10_932 ();
 FILLCELL_X2 FILLER_10_936 ();
 FILLCELL_X4 FILLER_10_945 ();
 FILLCELL_X2 FILLER_10_949 ();
 FILLCELL_X1 FILLER_10_953 ();
 FILLCELL_X8 FILLER_10_958 ();
 FILLCELL_X2 FILLER_10_966 ();
 FILLCELL_X4 FILLER_10_971 ();
 FILLCELL_X8 FILLER_10_997 ();
 FILLCELL_X1 FILLER_10_1005 ();
 FILLCELL_X2 FILLER_10_1028 ();
 FILLCELL_X8 FILLER_10_1035 ();
 FILLCELL_X1 FILLER_10_1052 ();
 FILLCELL_X1 FILLER_10_1058 ();
 FILLCELL_X1 FILLER_10_1068 ();
 FILLCELL_X2 FILLER_10_1091 ();
 FILLCELL_X1 FILLER_10_1093 ();
 FILLCELL_X1 FILLER_10_1114 ();
 FILLCELL_X8 FILLER_10_1122 ();
 FILLCELL_X1 FILLER_10_1135 ();
 FILLCELL_X1 FILLER_10_1209 ();
 FILLCELL_X16 FILLER_10_1237 ();
 FILLCELL_X2 FILLER_10_1253 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X16 FILLER_11_353 ();
 FILLCELL_X1 FILLER_11_369 ();
 FILLCELL_X2 FILLER_11_387 ();
 FILLCELL_X4 FILLER_11_406 ();
 FILLCELL_X1 FILLER_11_410 ();
 FILLCELL_X8 FILLER_11_442 ();
 FILLCELL_X1 FILLER_11_450 ();
 FILLCELL_X4 FILLER_11_460 ();
 FILLCELL_X2 FILLER_11_523 ();
 FILLCELL_X1 FILLER_11_525 ();
 FILLCELL_X2 FILLER_11_530 ();
 FILLCELL_X4 FILLER_11_541 ();
 FILLCELL_X2 FILLER_11_545 ();
 FILLCELL_X1 FILLER_11_547 ();
 FILLCELL_X8 FILLER_11_577 ();
 FILLCELL_X2 FILLER_11_585 ();
 FILLCELL_X2 FILLER_11_594 ();
 FILLCELL_X1 FILLER_11_596 ();
 FILLCELL_X2 FILLER_11_614 ();
 FILLCELL_X1 FILLER_11_616 ();
 FILLCELL_X4 FILLER_11_626 ();
 FILLCELL_X1 FILLER_11_630 ();
 FILLCELL_X4 FILLER_11_644 ();
 FILLCELL_X1 FILLER_11_648 ();
 FILLCELL_X4 FILLER_11_656 ();
 FILLCELL_X16 FILLER_11_667 ();
 FILLCELL_X4 FILLER_11_683 ();
 FILLCELL_X4 FILLER_11_707 ();
 FILLCELL_X2 FILLER_11_711 ();
 FILLCELL_X2 FILLER_11_718 ();
 FILLCELL_X2 FILLER_11_725 ();
 FILLCELL_X1 FILLER_11_734 ();
 FILLCELL_X1 FILLER_11_739 ();
 FILLCELL_X2 FILLER_11_743 ();
 FILLCELL_X1 FILLER_11_757 ();
 FILLCELL_X4 FILLER_11_767 ();
 FILLCELL_X1 FILLER_11_771 ();
 FILLCELL_X2 FILLER_11_776 ();
 FILLCELL_X1 FILLER_11_778 ();
 FILLCELL_X8 FILLER_11_806 ();
 FILLCELL_X4 FILLER_11_814 ();
 FILLCELL_X8 FILLER_11_828 ();
 FILLCELL_X1 FILLER_11_836 ();
 FILLCELL_X2 FILLER_11_842 ();
 FILLCELL_X1 FILLER_11_856 ();
 FILLCELL_X4 FILLER_11_864 ();
 FILLCELL_X1 FILLER_11_868 ();
 FILLCELL_X4 FILLER_11_886 ();
 FILLCELL_X2 FILLER_11_890 ();
 FILLCELL_X1 FILLER_11_901 ();
 FILLCELL_X2 FILLER_11_911 ();
 FILLCELL_X16 FILLER_11_920 ();
 FILLCELL_X1 FILLER_11_936 ();
 FILLCELL_X2 FILLER_11_942 ();
 FILLCELL_X2 FILLER_11_964 ();
 FILLCELL_X1 FILLER_11_966 ();
 FILLCELL_X1 FILLER_11_972 ();
 FILLCELL_X8 FILLER_11_988 ();
 FILLCELL_X4 FILLER_11_996 ();
 FILLCELL_X2 FILLER_11_1000 ();
 FILLCELL_X1 FILLER_11_1002 ();
 FILLCELL_X2 FILLER_11_1007 ();
 FILLCELL_X8 FILLER_11_1024 ();
 FILLCELL_X2 FILLER_11_1032 ();
 FILLCELL_X1 FILLER_11_1034 ();
 FILLCELL_X1 FILLER_11_1042 ();
 FILLCELL_X2 FILLER_11_1051 ();
 FILLCELL_X1 FILLER_11_1061 ();
 FILLCELL_X1 FILLER_11_1084 ();
 FILLCELL_X1 FILLER_11_1105 ();
 FILLCELL_X1 FILLER_11_1109 ();
 FILLCELL_X8 FILLER_11_1130 ();
 FILLCELL_X2 FILLER_11_1145 ();
 FILLCELL_X1 FILLER_11_1147 ();
 FILLCELL_X4 FILLER_11_1197 ();
 FILLCELL_X2 FILLER_11_1201 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X16 FILLER_12_353 ();
 FILLCELL_X4 FILLER_12_369 ();
 FILLCELL_X2 FILLER_12_373 ();
 FILLCELL_X1 FILLER_12_375 ();
 FILLCELL_X16 FILLER_12_397 ();
 FILLCELL_X4 FILLER_12_413 ();
 FILLCELL_X2 FILLER_12_417 ();
 FILLCELL_X16 FILLER_12_430 ();
 FILLCELL_X2 FILLER_12_446 ();
 FILLCELL_X4 FILLER_12_457 ();
 FILLCELL_X2 FILLER_12_461 ();
 FILLCELL_X1 FILLER_12_463 ();
 FILLCELL_X4 FILLER_12_481 ();
 FILLCELL_X2 FILLER_12_485 ();
 FILLCELL_X1 FILLER_12_487 ();
 FILLCELL_X8 FILLER_12_495 ();
 FILLCELL_X4 FILLER_12_503 ();
 FILLCELL_X2 FILLER_12_507 ();
 FILLCELL_X1 FILLER_12_509 ();
 FILLCELL_X2 FILLER_12_520 ();
 FILLCELL_X1 FILLER_12_522 ();
 FILLCELL_X2 FILLER_12_534 ();
 FILLCELL_X2 FILLER_12_545 ();
 FILLCELL_X1 FILLER_12_547 ();
 FILLCELL_X2 FILLER_12_552 ();
 FILLCELL_X2 FILLER_12_563 ();
 FILLCELL_X16 FILLER_12_572 ();
 FILLCELL_X2 FILLER_12_588 ();
 FILLCELL_X4 FILLER_12_595 ();
 FILLCELL_X2 FILLER_12_599 ();
 FILLCELL_X1 FILLER_12_601 ();
 FILLCELL_X1 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_617 ();
 FILLCELL_X2 FILLER_12_621 ();
 FILLCELL_X1 FILLER_12_623 ();
 FILLCELL_X2 FILLER_12_649 ();
 FILLCELL_X16 FILLER_12_675 ();
 FILLCELL_X4 FILLER_12_691 ();
 FILLCELL_X1 FILLER_12_739 ();
 FILLCELL_X2 FILLER_12_756 ();
 FILLCELL_X1 FILLER_12_758 ();
 FILLCELL_X2 FILLER_12_775 ();
 FILLCELL_X8 FILLER_12_822 ();
 FILLCELL_X4 FILLER_12_830 ();
 FILLCELL_X2 FILLER_12_834 ();
 FILLCELL_X1 FILLER_12_843 ();
 FILLCELL_X1 FILLER_12_848 ();
 FILLCELL_X1 FILLER_12_852 ();
 FILLCELL_X4 FILLER_12_877 ();
 FILLCELL_X1 FILLER_12_881 ();
 FILLCELL_X4 FILLER_12_925 ();
 FILLCELL_X1 FILLER_12_929 ();
 FILLCELL_X4 FILLER_12_945 ();
 FILLCELL_X1 FILLER_12_973 ();
 FILLCELL_X8 FILLER_12_978 ();
 FILLCELL_X4 FILLER_12_986 ();
 FILLCELL_X1 FILLER_12_990 ();
 FILLCELL_X1 FILLER_12_994 ();
 FILLCELL_X1 FILLER_12_999 ();
 FILLCELL_X2 FILLER_12_1007 ();
 FILLCELL_X1 FILLER_12_1016 ();
 FILLCELL_X2 FILLER_12_1021 ();
 FILLCELL_X1 FILLER_12_1023 ();
 FILLCELL_X4 FILLER_12_1032 ();
 FILLCELL_X2 FILLER_12_1036 ();
 FILLCELL_X4 FILLER_12_1041 ();
 FILLCELL_X8 FILLER_12_1082 ();
 FILLCELL_X4 FILLER_12_1090 ();
 FILLCELL_X4 FILLER_12_1147 ();
 FILLCELL_X2 FILLER_12_1151 ();
 FILLCELL_X4 FILLER_12_1167 ();
 FILLCELL_X2 FILLER_12_1175 ();
 FILLCELL_X2 FILLER_12_1180 ();
 FILLCELL_X2 FILLER_12_1202 ();
 FILLCELL_X2 FILLER_12_1211 ();
 FILLCELL_X32 FILLER_12_1220 ();
 FILLCELL_X2 FILLER_12_1252 ();
 FILLCELL_X1 FILLER_12_1254 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X16 FILLER_13_353 ();
 FILLCELL_X4 FILLER_13_369 ();
 FILLCELL_X2 FILLER_13_373 ();
 FILLCELL_X16 FILLER_13_382 ();
 FILLCELL_X4 FILLER_13_398 ();
 FILLCELL_X1 FILLER_13_402 ();
 FILLCELL_X1 FILLER_13_414 ();
 FILLCELL_X1 FILLER_13_422 ();
 FILLCELL_X16 FILLER_13_442 ();
 FILLCELL_X8 FILLER_13_458 ();
 FILLCELL_X2 FILLER_13_466 ();
 FILLCELL_X1 FILLER_13_471 ();
 FILLCELL_X8 FILLER_13_479 ();
 FILLCELL_X2 FILLER_13_487 ();
 FILLCELL_X2 FILLER_13_493 ();
 FILLCELL_X2 FILLER_13_511 ();
 FILLCELL_X2 FILLER_13_522 ();
 FILLCELL_X1 FILLER_13_524 ();
 FILLCELL_X4 FILLER_13_530 ();
 FILLCELL_X2 FILLER_13_545 ();
 FILLCELL_X1 FILLER_13_547 ();
 FILLCELL_X4 FILLER_13_561 ();
 FILLCELL_X1 FILLER_13_565 ();
 FILLCELL_X16 FILLER_13_571 ();
 FILLCELL_X4 FILLER_13_587 ();
 FILLCELL_X1 FILLER_13_603 ();
 FILLCELL_X8 FILLER_13_621 ();
 FILLCELL_X1 FILLER_13_629 ();
 FILLCELL_X2 FILLER_13_641 ();
 FILLCELL_X1 FILLER_13_643 ();
 FILLCELL_X2 FILLER_13_649 ();
 FILLCELL_X16 FILLER_13_667 ();
 FILLCELL_X4 FILLER_13_683 ();
 FILLCELL_X2 FILLER_13_687 ();
 FILLCELL_X1 FILLER_13_713 ();
 FILLCELL_X2 FILLER_13_717 ();
 FILLCELL_X2 FILLER_13_722 ();
 FILLCELL_X8 FILLER_13_726 ();
 FILLCELL_X2 FILLER_13_734 ();
 FILLCELL_X1 FILLER_13_736 ();
 FILLCELL_X16 FILLER_13_750 ();
 FILLCELL_X8 FILLER_13_766 ();
 FILLCELL_X4 FILLER_13_777 ();
 FILLCELL_X1 FILLER_13_781 ();
 FILLCELL_X2 FILLER_13_785 ();
 FILLCELL_X8 FILLER_13_808 ();
 FILLCELL_X2 FILLER_13_816 ();
 FILLCELL_X1 FILLER_13_818 ();
 FILLCELL_X2 FILLER_13_852 ();
 FILLCELL_X4 FILLER_13_861 ();
 FILLCELL_X4 FILLER_13_889 ();
 FILLCELL_X2 FILLER_13_893 ();
 FILLCELL_X4 FILLER_13_904 ();
 FILLCELL_X16 FILLER_13_915 ();
 FILLCELL_X4 FILLER_13_938 ();
 FILLCELL_X1 FILLER_13_942 ();
 FILLCELL_X2 FILLER_13_963 ();
 FILLCELL_X4 FILLER_13_995 ();
 FILLCELL_X1 FILLER_13_1004 ();
 FILLCELL_X1 FILLER_13_1009 ();
 FILLCELL_X2 FILLER_13_1018 ();
 FILLCELL_X1 FILLER_13_1020 ();
 FILLCELL_X4 FILLER_13_1025 ();
 FILLCELL_X1 FILLER_13_1029 ();
 FILLCELL_X2 FILLER_13_1034 ();
 FILLCELL_X1 FILLER_13_1036 ();
 FILLCELL_X2 FILLER_13_1050 ();
 FILLCELL_X16 FILLER_13_1061 ();
 FILLCELL_X8 FILLER_13_1077 ();
 FILLCELL_X2 FILLER_13_1085 ();
 FILLCELL_X1 FILLER_13_1117 ();
 FILLCELL_X2 FILLER_13_1123 ();
 FILLCELL_X16 FILLER_13_1145 ();
 FILLCELL_X8 FILLER_13_1161 ();
 FILLCELL_X2 FILLER_13_1169 ();
 FILLCELL_X4 FILLER_13_1193 ();
 FILLCELL_X1 FILLER_13_1197 ();
 FILLCELL_X16 FILLER_13_1238 ();
 FILLCELL_X1 FILLER_13_1254 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X8 FILLER_14_353 ();
 FILLCELL_X2 FILLER_14_361 ();
 FILLCELL_X1 FILLER_14_363 ();
 FILLCELL_X4 FILLER_14_381 ();
 FILLCELL_X2 FILLER_14_416 ();
 FILLCELL_X1 FILLER_14_418 ();
 FILLCELL_X4 FILLER_14_438 ();
 FILLCELL_X2 FILLER_14_442 ();
 FILLCELL_X1 FILLER_14_444 ();
 FILLCELL_X4 FILLER_14_485 ();
 FILLCELL_X1 FILLER_14_489 ();
 FILLCELL_X16 FILLER_14_510 ();
 FILLCELL_X8 FILLER_14_526 ();
 FILLCELL_X4 FILLER_14_534 ();
 FILLCELL_X8 FILLER_14_543 ();
 FILLCELL_X2 FILLER_14_551 ();
 FILLCELL_X1 FILLER_14_553 ();
 FILLCELL_X8 FILLER_14_572 ();
 FILLCELL_X1 FILLER_14_580 ();
 FILLCELL_X2 FILLER_14_590 ();
 FILLCELL_X4 FILLER_14_594 ();
 FILLCELL_X2 FILLER_14_598 ();
 FILLCELL_X8 FILLER_14_604 ();
 FILLCELL_X2 FILLER_14_612 ();
 FILLCELL_X2 FILLER_14_621 ();
 FILLCELL_X1 FILLER_14_623 ();
 FILLCELL_X1 FILLER_14_651 ();
 FILLCELL_X32 FILLER_14_659 ();
 FILLCELL_X4 FILLER_14_721 ();
 FILLCELL_X2 FILLER_14_725 ();
 FILLCELL_X1 FILLER_14_727 ();
 FILLCELL_X4 FILLER_14_730 ();
 FILLCELL_X2 FILLER_14_734 ();
 FILLCELL_X8 FILLER_14_740 ();
 FILLCELL_X4 FILLER_14_748 ();
 FILLCELL_X2 FILLER_14_752 ();
 FILLCELL_X4 FILLER_14_769 ();
 FILLCELL_X1 FILLER_14_773 ();
 FILLCELL_X2 FILLER_14_801 ();
 FILLCELL_X1 FILLER_14_803 ();
 FILLCELL_X2 FILLER_14_808 ();
 FILLCELL_X2 FILLER_14_817 ();
 FILLCELL_X1 FILLER_14_819 ();
 FILLCELL_X2 FILLER_14_825 ();
 FILLCELL_X1 FILLER_14_827 ();
 FILLCELL_X2 FILLER_14_831 ();
 FILLCELL_X1 FILLER_14_833 ();
 FILLCELL_X2 FILLER_14_845 ();
 FILLCELL_X8 FILLER_14_854 ();
 FILLCELL_X1 FILLER_14_862 ();
 FILLCELL_X16 FILLER_14_876 ();
 FILLCELL_X4 FILLER_14_892 ();
 FILLCELL_X2 FILLER_14_896 ();
 FILLCELL_X4 FILLER_14_907 ();
 FILLCELL_X4 FILLER_14_941 ();
 FILLCELL_X2 FILLER_14_945 ();
 FILLCELL_X4 FILLER_14_950 ();
 FILLCELL_X2 FILLER_14_954 ();
 FILLCELL_X1 FILLER_14_956 ();
 FILLCELL_X2 FILLER_14_979 ();
 FILLCELL_X4 FILLER_14_988 ();
 FILLCELL_X1 FILLER_14_992 ();
 FILLCELL_X2 FILLER_14_1020 ();
 FILLCELL_X8 FILLER_14_1026 ();
 FILLCELL_X2 FILLER_14_1034 ();
 FILLCELL_X1 FILLER_14_1036 ();
 FILLCELL_X4 FILLER_14_1059 ();
 FILLCELL_X2 FILLER_14_1063 ();
 FILLCELL_X1 FILLER_14_1065 ();
 FILLCELL_X4 FILLER_14_1088 ();
 FILLCELL_X1 FILLER_14_1092 ();
 FILLCELL_X2 FILLER_14_1100 ();
 FILLCELL_X1 FILLER_14_1107 ();
 FILLCELL_X4 FILLER_14_1135 ();
 FILLCELL_X8 FILLER_14_1146 ();
 FILLCELL_X1 FILLER_14_1154 ();
 FILLCELL_X1 FILLER_14_1184 ();
 FILLCELL_X8 FILLER_14_1210 ();
 FILLCELL_X2 FILLER_14_1218 ();
 FILLCELL_X1 FILLER_14_1220 ();
 FILLCELL_X4 FILLER_14_1250 ();
 FILLCELL_X1 FILLER_14_1254 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X16 FILLER_15_353 ();
 FILLCELL_X8 FILLER_15_369 ();
 FILLCELL_X2 FILLER_15_377 ();
 FILLCELL_X1 FILLER_15_379 ();
 FILLCELL_X1 FILLER_15_387 ();
 FILLCELL_X2 FILLER_15_393 ();
 FILLCELL_X8 FILLER_15_419 ();
 FILLCELL_X1 FILLER_15_427 ();
 FILLCELL_X1 FILLER_15_445 ();
 FILLCELL_X1 FILLER_15_453 ();
 FILLCELL_X1 FILLER_15_458 ();
 FILLCELL_X4 FILLER_15_489 ();
 FILLCELL_X1 FILLER_15_502 ();
 FILLCELL_X2 FILLER_15_512 ();
 FILLCELL_X2 FILLER_15_519 ();
 FILLCELL_X2 FILLER_15_526 ();
 FILLCELL_X1 FILLER_15_533 ();
 FILLCELL_X2 FILLER_15_549 ();
 FILLCELL_X1 FILLER_15_562 ();
 FILLCELL_X2 FILLER_15_571 ();
 FILLCELL_X2 FILLER_15_577 ();
 FILLCELL_X1 FILLER_15_586 ();
 FILLCELL_X8 FILLER_15_596 ();
 FILLCELL_X1 FILLER_15_604 ();
 FILLCELL_X4 FILLER_15_614 ();
 FILLCELL_X8 FILLER_15_625 ();
 FILLCELL_X8 FILLER_15_646 ();
 FILLCELL_X1 FILLER_15_671 ();
 FILLCELL_X4 FILLER_15_696 ();
 FILLCELL_X1 FILLER_15_700 ();
 FILLCELL_X4 FILLER_15_705 ();
 FILLCELL_X1 FILLER_15_731 ();
 FILLCELL_X1 FILLER_15_742 ();
 FILLCELL_X1 FILLER_15_748 ();
 FILLCELL_X1 FILLER_15_771 ();
 FILLCELL_X4 FILLER_15_778 ();
 FILLCELL_X1 FILLER_15_782 ();
 FILLCELL_X1 FILLER_15_791 ();
 FILLCELL_X2 FILLER_15_829 ();
 FILLCELL_X1 FILLER_15_839 ();
 FILLCELL_X1 FILLER_15_854 ();
 FILLCELL_X4 FILLER_15_859 ();
 FILLCELL_X2 FILLER_15_863 ();
 FILLCELL_X16 FILLER_15_868 ();
 FILLCELL_X2 FILLER_15_884 ();
 FILLCELL_X2 FILLER_15_893 ();
 FILLCELL_X4 FILLER_15_900 ();
 FILLCELL_X1 FILLER_15_904 ();
 FILLCELL_X8 FILLER_15_927 ();
 FILLCELL_X4 FILLER_15_939 ();
 FILLCELL_X1 FILLER_15_943 ();
 FILLCELL_X4 FILLER_15_948 ();
 FILLCELL_X2 FILLER_15_970 ();
 FILLCELL_X1 FILLER_15_985 ();
 FILLCELL_X4 FILLER_15_1006 ();
 FILLCELL_X2 FILLER_15_1010 ();
 FILLCELL_X1 FILLER_15_1012 ();
 FILLCELL_X16 FILLER_15_1033 ();
 FILLCELL_X8 FILLER_15_1049 ();
 FILLCELL_X4 FILLER_15_1057 ();
 FILLCELL_X1 FILLER_15_1079 ();
 FILLCELL_X4 FILLER_15_1109 ();
 FILLCELL_X1 FILLER_15_1113 ();
 FILLCELL_X8 FILLER_15_1126 ();
 FILLCELL_X4 FILLER_15_1134 ();
 FILLCELL_X16 FILLER_15_1160 ();
 FILLCELL_X2 FILLER_15_1183 ();
 FILLCELL_X1 FILLER_15_1189 ();
 FILLCELL_X4 FILLER_15_1194 ();
 FILLCELL_X16 FILLER_15_1236 ();
 FILLCELL_X2 FILLER_15_1252 ();
 FILLCELL_X1 FILLER_15_1254 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X16 FILLER_16_353 ();
 FILLCELL_X4 FILLER_16_369 ();
 FILLCELL_X2 FILLER_16_373 ();
 FILLCELL_X1 FILLER_16_375 ();
 FILLCELL_X2 FILLER_16_383 ();
 FILLCELL_X2 FILLER_16_426 ();
 FILLCELL_X1 FILLER_16_428 ();
 FILLCELL_X1 FILLER_16_439 ();
 FILLCELL_X1 FILLER_16_447 ();
 FILLCELL_X1 FILLER_16_455 ();
 FILLCELL_X1 FILLER_16_469 ();
 FILLCELL_X8 FILLER_16_484 ();
 FILLCELL_X1 FILLER_16_503 ();
 FILLCELL_X2 FILLER_16_515 ();
 FILLCELL_X2 FILLER_16_521 ();
 FILLCELL_X1 FILLER_16_523 ();
 FILLCELL_X1 FILLER_16_550 ();
 FILLCELL_X1 FILLER_16_576 ();
 FILLCELL_X1 FILLER_16_581 ();
 FILLCELL_X2 FILLER_16_590 ();
 FILLCELL_X1 FILLER_16_597 ();
 FILLCELL_X4 FILLER_16_602 ();
 FILLCELL_X4 FILLER_16_611 ();
 FILLCELL_X2 FILLER_16_615 ();
 FILLCELL_X1 FILLER_16_621 ();
 FILLCELL_X8 FILLER_16_643 ();
 FILLCELL_X8 FILLER_16_664 ();
 FILLCELL_X4 FILLER_16_672 ();
 FILLCELL_X2 FILLER_16_676 ();
 FILLCELL_X4 FILLER_16_698 ();
 FILLCELL_X1 FILLER_16_702 ();
 FILLCELL_X1 FILLER_16_707 ();
 FILLCELL_X1 FILLER_16_728 ();
 FILLCELL_X1 FILLER_16_733 ();
 FILLCELL_X4 FILLER_16_747 ();
 FILLCELL_X1 FILLER_16_751 ();
 FILLCELL_X2 FILLER_16_756 ();
 FILLCELL_X2 FILLER_16_762 ();
 FILLCELL_X1 FILLER_16_764 ();
 FILLCELL_X1 FILLER_16_770 ();
 FILLCELL_X2 FILLER_16_778 ();
 FILLCELL_X1 FILLER_16_780 ();
 FILLCELL_X16 FILLER_16_807 ();
 FILLCELL_X4 FILLER_16_823 ();
 FILLCELL_X2 FILLER_16_827 ();
 FILLCELL_X1 FILLER_16_829 ();
 FILLCELL_X4 FILLER_16_840 ();
 FILLCELL_X2 FILLER_16_855 ();
 FILLCELL_X8 FILLER_16_879 ();
 FILLCELL_X4 FILLER_16_887 ();
 FILLCELL_X1 FILLER_16_891 ();
 FILLCELL_X2 FILLER_16_927 ();
 FILLCELL_X2 FILLER_16_931 ();
 FILLCELL_X1 FILLER_16_951 ();
 FILLCELL_X4 FILLER_16_956 ();
 FILLCELL_X2 FILLER_16_960 ();
 FILLCELL_X8 FILLER_16_965 ();
 FILLCELL_X2 FILLER_16_976 ();
 FILLCELL_X8 FILLER_16_1010 ();
 FILLCELL_X4 FILLER_16_1023 ();
 FILLCELL_X1 FILLER_16_1027 ();
 FILLCELL_X2 FILLER_16_1059 ();
 FILLCELL_X8 FILLER_16_1068 ();
 FILLCELL_X1 FILLER_16_1076 ();
 FILLCELL_X8 FILLER_16_1097 ();
 FILLCELL_X1 FILLER_16_1105 ();
 FILLCELL_X4 FILLER_16_1109 ();
 FILLCELL_X8 FILLER_16_1147 ();
 FILLCELL_X1 FILLER_16_1155 ();
 FILLCELL_X2 FILLER_16_1181 ();
 FILLCELL_X4 FILLER_16_1205 ();
 FILLCELL_X2 FILLER_16_1209 ();
 FILLCELL_X4 FILLER_16_1216 ();
 FILLCELL_X2 FILLER_16_1222 ();
 FILLCELL_X1 FILLER_16_1224 ();
 FILLCELL_X4 FILLER_16_1250 ();
 FILLCELL_X1 FILLER_16_1254 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X8 FILLER_17_353 ();
 FILLCELL_X2 FILLER_17_361 ();
 FILLCELL_X1 FILLER_17_363 ();
 FILLCELL_X2 FILLER_17_381 ();
 FILLCELL_X16 FILLER_17_390 ();
 FILLCELL_X8 FILLER_17_406 ();
 FILLCELL_X4 FILLER_17_414 ();
 FILLCELL_X1 FILLER_17_418 ();
 FILLCELL_X2 FILLER_17_433 ();
 FILLCELL_X16 FILLER_17_440 ();
 FILLCELL_X1 FILLER_17_456 ();
 FILLCELL_X32 FILLER_17_461 ();
 FILLCELL_X4 FILLER_17_497 ();
 FILLCELL_X2 FILLER_17_501 ();
 FILLCELL_X2 FILLER_17_507 ();
 FILLCELL_X1 FILLER_17_516 ();
 FILLCELL_X1 FILLER_17_521 ();
 FILLCELL_X4 FILLER_17_530 ();
 FILLCELL_X2 FILLER_17_534 ();
 FILLCELL_X2 FILLER_17_558 ();
 FILLCELL_X2 FILLER_17_567 ();
 FILLCELL_X1 FILLER_17_569 ();
 FILLCELL_X2 FILLER_17_577 ();
 FILLCELL_X2 FILLER_17_611 ();
 FILLCELL_X4 FILLER_17_628 ();
 FILLCELL_X2 FILLER_17_632 ();
 FILLCELL_X4 FILLER_17_647 ();
 FILLCELL_X1 FILLER_17_651 ();
 FILLCELL_X1 FILLER_17_654 ();
 FILLCELL_X8 FILLER_17_659 ();
 FILLCELL_X8 FILLER_17_678 ();
 FILLCELL_X4 FILLER_17_686 ();
 FILLCELL_X4 FILLER_17_712 ();
 FILLCELL_X16 FILLER_17_727 ();
 FILLCELL_X4 FILLER_17_743 ();
 FILLCELL_X2 FILLER_17_759 ();
 FILLCELL_X1 FILLER_17_761 ();
 FILLCELL_X16 FILLER_17_777 ();
 FILLCELL_X4 FILLER_17_793 ();
 FILLCELL_X2 FILLER_17_797 ();
 FILLCELL_X2 FILLER_17_803 ();
 FILLCELL_X1 FILLER_17_805 ();
 FILLCELL_X1 FILLER_17_839 ();
 FILLCELL_X2 FILLER_17_848 ();
 FILLCELL_X8 FILLER_17_854 ();
 FILLCELL_X1 FILLER_17_862 ();
 FILLCELL_X2 FILLER_17_885 ();
 FILLCELL_X4 FILLER_17_905 ();
 FILLCELL_X2 FILLER_17_909 ();
 FILLCELL_X1 FILLER_17_911 ();
 FILLCELL_X2 FILLER_17_917 ();
 FILLCELL_X2 FILLER_17_934 ();
 FILLCELL_X4 FILLER_17_945 ();
 FILLCELL_X2 FILLER_17_949 ();
 FILLCELL_X1 FILLER_17_954 ();
 FILLCELL_X2 FILLER_17_958 ();
 FILLCELL_X2 FILLER_17_988 ();
 FILLCELL_X8 FILLER_17_997 ();
 FILLCELL_X1 FILLER_17_1005 ();
 FILLCELL_X4 FILLER_17_1033 ();
 FILLCELL_X1 FILLER_17_1037 ();
 FILLCELL_X4 FILLER_17_1078 ();
 FILLCELL_X1 FILLER_17_1082 ();
 FILLCELL_X4 FILLER_17_1094 ();
 FILLCELL_X1 FILLER_17_1098 ();
 FILLCELL_X4 FILLER_17_1106 ();
 FILLCELL_X2 FILLER_17_1110 ();
 FILLCELL_X4 FILLER_17_1119 ();
 FILLCELL_X4 FILLER_17_1132 ();
 FILLCELL_X2 FILLER_17_1136 ();
 FILLCELL_X4 FILLER_17_1167 ();
 FILLCELL_X2 FILLER_17_1171 ();
 FILLCELL_X1 FILLER_17_1173 ();
 FILLCELL_X2 FILLER_17_1185 ();
 FILLCELL_X4 FILLER_17_1190 ();
 FILLCELL_X4 FILLER_17_1201 ();
 FILLCELL_X2 FILLER_17_1205 ();
 FILLCELL_X1 FILLER_17_1207 ();
 FILLCELL_X1 FILLER_17_1213 ();
 FILLCELL_X4 FILLER_17_1221 ();
 FILLCELL_X1 FILLER_17_1225 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X16 FILLER_18_353 ();
 FILLCELL_X8 FILLER_18_369 ();
 FILLCELL_X2 FILLER_18_377 ();
 FILLCELL_X4 FILLER_18_386 ();
 FILLCELL_X1 FILLER_18_390 ();
 FILLCELL_X4 FILLER_18_415 ();
 FILLCELL_X2 FILLER_18_443 ();
 FILLCELL_X1 FILLER_18_445 ();
 FILLCELL_X2 FILLER_18_455 ();
 FILLCELL_X2 FILLER_18_464 ();
 FILLCELL_X2 FILLER_18_470 ();
 FILLCELL_X4 FILLER_18_485 ();
 FILLCELL_X1 FILLER_18_489 ();
 FILLCELL_X4 FILLER_18_497 ();
 FILLCELL_X1 FILLER_18_501 ();
 FILLCELL_X1 FILLER_18_519 ();
 FILLCELL_X16 FILLER_18_543 ();
 FILLCELL_X2 FILLER_18_571 ();
 FILLCELL_X1 FILLER_18_573 ();
 FILLCELL_X2 FILLER_18_607 ();
 FILLCELL_X1 FILLER_18_609 ();
 FILLCELL_X8 FILLER_18_621 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X2 FILLER_18_648 ();
 FILLCELL_X1 FILLER_18_650 ();
 FILLCELL_X8 FILLER_18_659 ();
 FILLCELL_X1 FILLER_18_671 ();
 FILLCELL_X4 FILLER_18_680 ();
 FILLCELL_X1 FILLER_18_692 ();
 FILLCELL_X2 FILLER_18_721 ();
 FILLCELL_X1 FILLER_18_759 ();
 FILLCELL_X2 FILLER_18_793 ();
 FILLCELL_X1 FILLER_18_795 ();
 FILLCELL_X8 FILLER_18_825 ();
 FILLCELL_X16 FILLER_18_870 ();
 FILLCELL_X2 FILLER_18_886 ();
 FILLCELL_X1 FILLER_18_908 ();
 FILLCELL_X1 FILLER_18_912 ();
 FILLCELL_X1 FILLER_18_926 ();
 FILLCELL_X8 FILLER_18_939 ();
 FILLCELL_X1 FILLER_18_947 ();
 FILLCELL_X16 FILLER_18_955 ();
 FILLCELL_X16 FILLER_18_1009 ();
 FILLCELL_X8 FILLER_18_1025 ();
 FILLCELL_X4 FILLER_18_1033 ();
 FILLCELL_X2 FILLER_18_1037 ();
 FILLCELL_X4 FILLER_18_1053 ();
 FILLCELL_X2 FILLER_18_1057 ();
 FILLCELL_X8 FILLER_18_1066 ();
 FILLCELL_X2 FILLER_18_1074 ();
 FILLCELL_X1 FILLER_18_1076 ();
 FILLCELL_X2 FILLER_18_1129 ();
 FILLCELL_X1 FILLER_18_1143 ();
 FILLCELL_X1 FILLER_18_1151 ();
 FILLCELL_X1 FILLER_18_1189 ();
 FILLCELL_X2 FILLER_18_1210 ();
 FILLCELL_X1 FILLER_18_1212 ();
 FILLCELL_X2 FILLER_18_1233 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X16 FILLER_19_353 ();
 FILLCELL_X4 FILLER_19_369 ();
 FILLCELL_X4 FILLER_19_397 ();
 FILLCELL_X1 FILLER_19_401 ();
 FILLCELL_X4 FILLER_19_419 ();
 FILLCELL_X8 FILLER_19_460 ();
 FILLCELL_X1 FILLER_19_468 ();
 FILLCELL_X8 FILLER_19_478 ();
 FILLCELL_X2 FILLER_19_486 ();
 FILLCELL_X1 FILLER_19_488 ();
 FILLCELL_X4 FILLER_19_498 ();
 FILLCELL_X2 FILLER_19_502 ();
 FILLCELL_X2 FILLER_19_513 ();
 FILLCELL_X1 FILLER_19_530 ();
 FILLCELL_X2 FILLER_19_557 ();
 FILLCELL_X2 FILLER_19_563 ();
 FILLCELL_X2 FILLER_19_597 ();
 FILLCELL_X2 FILLER_19_624 ();
 FILLCELL_X1 FILLER_19_626 ();
 FILLCELL_X4 FILLER_19_634 ();
 FILLCELL_X1 FILLER_19_638 ();
 FILLCELL_X8 FILLER_19_646 ();
 FILLCELL_X4 FILLER_19_654 ();
 FILLCELL_X2 FILLER_19_658 ();
 FILLCELL_X4 FILLER_19_664 ();
 FILLCELL_X8 FILLER_19_672 ();
 FILLCELL_X1 FILLER_19_680 ();
 FILLCELL_X2 FILLER_19_688 ();
 FILLCELL_X8 FILLER_19_710 ();
 FILLCELL_X2 FILLER_19_718 ();
 FILLCELL_X1 FILLER_19_720 ();
 FILLCELL_X2 FILLER_19_730 ();
 FILLCELL_X1 FILLER_19_737 ();
 FILLCELL_X2 FILLER_19_743 ();
 FILLCELL_X2 FILLER_19_748 ();
 FILLCELL_X2 FILLER_19_759 ();
 FILLCELL_X4 FILLER_19_764 ();
 FILLCELL_X1 FILLER_19_768 ();
 FILLCELL_X1 FILLER_19_780 ();
 FILLCELL_X2 FILLER_19_788 ();
 FILLCELL_X1 FILLER_19_790 ();
 FILLCELL_X2 FILLER_19_796 ();
 FILLCELL_X2 FILLER_19_812 ();
 FILLCELL_X1 FILLER_19_817 ();
 FILLCELL_X16 FILLER_19_835 ();
 FILLCELL_X1 FILLER_19_851 ();
 FILLCELL_X2 FILLER_19_855 ();
 FILLCELL_X1 FILLER_19_857 ();
 FILLCELL_X2 FILLER_19_864 ();
 FILLCELL_X1 FILLER_19_880 ();
 FILLCELL_X4 FILLER_19_890 ();
 FILLCELL_X2 FILLER_19_894 ();
 FILLCELL_X1 FILLER_19_896 ();
 FILLCELL_X2 FILLER_19_918 ();
 FILLCELL_X1 FILLER_19_920 ();
 FILLCELL_X4 FILLER_19_924 ();
 FILLCELL_X2 FILLER_19_969 ();
 FILLCELL_X1 FILLER_19_991 ();
 FILLCELL_X4 FILLER_19_1000 ();
 FILLCELL_X1 FILLER_19_1004 ();
 FILLCELL_X4 FILLER_19_1052 ();
 FILLCELL_X8 FILLER_19_1076 ();
 FILLCELL_X1 FILLER_19_1084 ();
 FILLCELL_X4 FILLER_19_1088 ();
 FILLCELL_X2 FILLER_19_1097 ();
 FILLCELL_X32 FILLER_19_1133 ();
 FILLCELL_X2 FILLER_19_1169 ();
 FILLCELL_X16 FILLER_19_1180 ();
 FILLCELL_X8 FILLER_19_1196 ();
 FILLCELL_X1 FILLER_19_1208 ();
 FILLCELL_X1 FILLER_19_1212 ();
 FILLCELL_X8 FILLER_19_1244 ();
 FILLCELL_X2 FILLER_19_1252 ();
 FILLCELL_X1 FILLER_19_1254 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X16 FILLER_20_392 ();
 FILLCELL_X2 FILLER_20_408 ();
 FILLCELL_X1 FILLER_20_417 ();
 FILLCELL_X1 FILLER_20_425 ();
 FILLCELL_X1 FILLER_20_433 ();
 FILLCELL_X4 FILLER_20_448 ();
 FILLCELL_X1 FILLER_20_452 ();
 FILLCELL_X2 FILLER_20_459 ();
 FILLCELL_X1 FILLER_20_461 ();
 FILLCELL_X2 FILLER_20_469 ();
 FILLCELL_X1 FILLER_20_478 ();
 FILLCELL_X1 FILLER_20_486 ();
 FILLCELL_X2 FILLER_20_492 ();
 FILLCELL_X4 FILLER_20_510 ();
 FILLCELL_X2 FILLER_20_514 ();
 FILLCELL_X4 FILLER_20_523 ();
 FILLCELL_X2 FILLER_20_527 ();
 FILLCELL_X1 FILLER_20_529 ();
 FILLCELL_X2 FILLER_20_541 ();
 FILLCELL_X1 FILLER_20_543 ();
 FILLCELL_X1 FILLER_20_549 ();
 FILLCELL_X2 FILLER_20_554 ();
 FILLCELL_X2 FILLER_20_560 ();
 FILLCELL_X1 FILLER_20_573 ();
 FILLCELL_X4 FILLER_20_580 ();
 FILLCELL_X1 FILLER_20_584 ();
 FILLCELL_X1 FILLER_20_593 ();
 FILLCELL_X1 FILLER_20_604 ();
 FILLCELL_X2 FILLER_20_620 ();
 FILLCELL_X4 FILLER_20_626 ();
 FILLCELL_X1 FILLER_20_630 ();
 FILLCELL_X8 FILLER_20_632 ();
 FILLCELL_X2 FILLER_20_640 ();
 FILLCELL_X16 FILLER_20_663 ();
 FILLCELL_X4 FILLER_20_699 ();
 FILLCELL_X1 FILLER_20_740 ();
 FILLCELL_X1 FILLER_20_745 ();
 FILLCELL_X4 FILLER_20_750 ();
 FILLCELL_X1 FILLER_20_754 ();
 FILLCELL_X8 FILLER_20_758 ();
 FILLCELL_X4 FILLER_20_766 ();
 FILLCELL_X2 FILLER_20_770 ();
 FILLCELL_X1 FILLER_20_772 ();
 FILLCELL_X1 FILLER_20_779 ();
 FILLCELL_X2 FILLER_20_788 ();
 FILLCELL_X2 FILLER_20_795 ();
 FILLCELL_X1 FILLER_20_797 ();
 FILLCELL_X1 FILLER_20_803 ();
 FILLCELL_X2 FILLER_20_807 ();
 FILLCELL_X2 FILLER_20_813 ();
 FILLCELL_X2 FILLER_20_819 ();
 FILLCELL_X2 FILLER_20_825 ();
 FILLCELL_X1 FILLER_20_827 ();
 FILLCELL_X2 FILLER_20_857 ();
 FILLCELL_X1 FILLER_20_867 ();
 FILLCELL_X2 FILLER_20_871 ();
 FILLCELL_X2 FILLER_20_878 ();
 FILLCELL_X1 FILLER_20_880 ();
 FILLCELL_X2 FILLER_20_886 ();
 FILLCELL_X8 FILLER_20_907 ();
 FILLCELL_X4 FILLER_20_925 ();
 FILLCELL_X1 FILLER_20_929 ();
 FILLCELL_X1 FILLER_20_934 ();
 FILLCELL_X1 FILLER_20_955 ();
 FILLCELL_X8 FILLER_20_974 ();
 FILLCELL_X1 FILLER_20_982 ();
 FILLCELL_X1 FILLER_20_987 ();
 FILLCELL_X8 FILLER_20_992 ();
 FILLCELL_X4 FILLER_20_1000 ();
 FILLCELL_X1 FILLER_20_1004 ();
 FILLCELL_X8 FILLER_20_1012 ();
 FILLCELL_X2 FILLER_20_1020 ();
 FILLCELL_X8 FILLER_20_1024 ();
 FILLCELL_X4 FILLER_20_1032 ();
 FILLCELL_X2 FILLER_20_1036 ();
 FILLCELL_X1 FILLER_20_1038 ();
 FILLCELL_X8 FILLER_20_1048 ();
 FILLCELL_X1 FILLER_20_1056 ();
 FILLCELL_X1 FILLER_20_1077 ();
 FILLCELL_X4 FILLER_20_1100 ();
 FILLCELL_X1 FILLER_20_1132 ();
 FILLCELL_X4 FILLER_20_1184 ();
 FILLCELL_X1 FILLER_20_1188 ();
 FILLCELL_X8 FILLER_20_1192 ();
 FILLCELL_X16 FILLER_20_1228 ();
 FILLCELL_X8 FILLER_20_1244 ();
 FILLCELL_X2 FILLER_20_1252 ();
 FILLCELL_X1 FILLER_20_1254 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X16 FILLER_21_353 ();
 FILLCELL_X4 FILLER_21_369 ();
 FILLCELL_X16 FILLER_21_387 ();
 FILLCELL_X4 FILLER_21_403 ();
 FILLCELL_X2 FILLER_21_414 ();
 FILLCELL_X1 FILLER_21_416 ();
 FILLCELL_X8 FILLER_21_422 ();
 FILLCELL_X2 FILLER_21_430 ();
 FILLCELL_X1 FILLER_21_432 ();
 FILLCELL_X2 FILLER_21_470 ();
 FILLCELL_X1 FILLER_21_472 ();
 FILLCELL_X16 FILLER_21_486 ();
 FILLCELL_X2 FILLER_21_502 ();
 FILLCELL_X1 FILLER_21_516 ();
 FILLCELL_X4 FILLER_21_527 ();
 FILLCELL_X1 FILLER_21_546 ();
 FILLCELL_X4 FILLER_21_555 ();
 FILLCELL_X1 FILLER_21_583 ();
 FILLCELL_X2 FILLER_21_592 ();
 FILLCELL_X2 FILLER_21_626 ();
 FILLCELL_X1 FILLER_21_633 ();
 FILLCELL_X4 FILLER_21_643 ();
 FILLCELL_X2 FILLER_21_647 ();
 FILLCELL_X2 FILLER_21_667 ();
 FILLCELL_X1 FILLER_21_669 ();
 FILLCELL_X16 FILLER_21_677 ();
 FILLCELL_X4 FILLER_21_693 ();
 FILLCELL_X1 FILLER_21_707 ();
 FILLCELL_X1 FILLER_21_711 ();
 FILLCELL_X1 FILLER_21_721 ();
 FILLCELL_X2 FILLER_21_745 ();
 FILLCELL_X1 FILLER_21_752 ();
 FILLCELL_X1 FILLER_21_757 ();
 FILLCELL_X1 FILLER_21_762 ();
 FILLCELL_X4 FILLER_21_774 ();
 FILLCELL_X2 FILLER_21_778 ();
 FILLCELL_X2 FILLER_21_785 ();
 FILLCELL_X1 FILLER_21_787 ();
 FILLCELL_X1 FILLER_21_821 ();
 FILLCELL_X1 FILLER_21_829 ();
 FILLCELL_X4 FILLER_21_852 ();
 FILLCELL_X2 FILLER_21_856 ();
 FILLCELL_X2 FILLER_21_908 ();
 FILLCELL_X8 FILLER_21_934 ();
 FILLCELL_X4 FILLER_21_942 ();
 FILLCELL_X1 FILLER_21_946 ();
 FILLCELL_X1 FILLER_21_968 ();
 FILLCELL_X8 FILLER_21_989 ();
 FILLCELL_X4 FILLER_21_1017 ();
 FILLCELL_X2 FILLER_21_1021 ();
 FILLCELL_X1 FILLER_21_1030 ();
 FILLCELL_X2 FILLER_21_1038 ();
 FILLCELL_X1 FILLER_21_1067 ();
 FILLCELL_X8 FILLER_21_1082 ();
 FILLCELL_X2 FILLER_21_1097 ();
 FILLCELL_X2 FILLER_21_1106 ();
 FILLCELL_X1 FILLER_21_1108 ();
 FILLCELL_X1 FILLER_21_1112 ();
 FILLCELL_X16 FILLER_21_1147 ();
 FILLCELL_X2 FILLER_21_1163 ();
 FILLCELL_X1 FILLER_21_1165 ();
 FILLCELL_X1 FILLER_21_1175 ();
 FILLCELL_X4 FILLER_21_1206 ();
 FILLCELL_X4 FILLER_21_1222 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X8 FILLER_22_353 ();
 FILLCELL_X4 FILLER_22_361 ();
 FILLCELL_X1 FILLER_22_365 ();
 FILLCELL_X1 FILLER_22_383 ();
 FILLCELL_X4 FILLER_22_391 ();
 FILLCELL_X2 FILLER_22_395 ();
 FILLCELL_X1 FILLER_22_397 ();
 FILLCELL_X16 FILLER_22_420 ();
 FILLCELL_X4 FILLER_22_436 ();
 FILLCELL_X2 FILLER_22_440 ();
 FILLCELL_X2 FILLER_22_449 ();
 FILLCELL_X1 FILLER_22_480 ();
 FILLCELL_X4 FILLER_22_490 ();
 FILLCELL_X2 FILLER_22_494 ();
 FILLCELL_X2 FILLER_22_513 ();
 FILLCELL_X8 FILLER_22_525 ();
 FILLCELL_X4 FILLER_22_539 ();
 FILLCELL_X2 FILLER_22_543 ();
 FILLCELL_X2 FILLER_22_563 ();
 FILLCELL_X1 FILLER_22_570 ();
 FILLCELL_X4 FILLER_22_582 ();
 FILLCELL_X2 FILLER_22_586 ();
 FILLCELL_X1 FILLER_22_588 ();
 FILLCELL_X4 FILLER_22_602 ();
 FILLCELL_X1 FILLER_22_606 ();
 FILLCELL_X1 FILLER_22_612 ();
 FILLCELL_X2 FILLER_22_620 ();
 FILLCELL_X4 FILLER_22_626 ();
 FILLCELL_X1 FILLER_22_630 ();
 FILLCELL_X8 FILLER_22_632 ();
 FILLCELL_X4 FILLER_22_640 ();
 FILLCELL_X2 FILLER_22_644 ();
 FILLCELL_X8 FILLER_22_653 ();
 FILLCELL_X4 FILLER_22_661 ();
 FILLCELL_X2 FILLER_22_672 ();
 FILLCELL_X1 FILLER_22_674 ();
 FILLCELL_X8 FILLER_22_680 ();
 FILLCELL_X4 FILLER_22_688 ();
 FILLCELL_X2 FILLER_22_692 ();
 FILLCELL_X1 FILLER_22_694 ();
 FILLCELL_X1 FILLER_22_702 ();
 FILLCELL_X1 FILLER_22_707 ();
 FILLCELL_X1 FILLER_22_712 ();
 FILLCELL_X1 FILLER_22_717 ();
 FILLCELL_X1 FILLER_22_722 ();
 FILLCELL_X1 FILLER_22_749 ();
 FILLCELL_X1 FILLER_22_754 ();
 FILLCELL_X1 FILLER_22_757 ();
 FILLCELL_X1 FILLER_22_761 ();
 FILLCELL_X8 FILLER_22_774 ();
 FILLCELL_X2 FILLER_22_782 ();
 FILLCELL_X1 FILLER_22_784 ();
 FILLCELL_X2 FILLER_22_795 ();
 FILLCELL_X2 FILLER_22_800 ();
 FILLCELL_X4 FILLER_22_817 ();
 FILLCELL_X2 FILLER_22_821 ();
 FILLCELL_X1 FILLER_22_823 ();
 FILLCELL_X8 FILLER_22_829 ();
 FILLCELL_X1 FILLER_22_837 ();
 FILLCELL_X8 FILLER_22_849 ();
 FILLCELL_X4 FILLER_22_857 ();
 FILLCELL_X1 FILLER_22_861 ();
 FILLCELL_X32 FILLER_22_867 ();
 FILLCELL_X2 FILLER_22_899 ();
 FILLCELL_X4 FILLER_22_912 ();
 FILLCELL_X2 FILLER_22_916 ();
 FILLCELL_X1 FILLER_22_918 ();
 FILLCELL_X8 FILLER_22_927 ();
 FILLCELL_X2 FILLER_22_935 ();
 FILLCELL_X1 FILLER_22_937 ();
 FILLCELL_X4 FILLER_22_952 ();
 FILLCELL_X2 FILLER_22_956 ();
 FILLCELL_X1 FILLER_22_958 ();
 FILLCELL_X2 FILLER_22_967 ();
 FILLCELL_X2 FILLER_22_973 ();
 FILLCELL_X2 FILLER_22_986 ();
 FILLCELL_X2 FILLER_22_1008 ();
 FILLCELL_X1 FILLER_22_1010 ();
 FILLCELL_X2 FILLER_22_1051 ();
 FILLCELL_X1 FILLER_22_1053 ();
 FILLCELL_X1 FILLER_22_1061 ();
 FILLCELL_X2 FILLER_22_1087 ();
 FILLCELL_X2 FILLER_22_1109 ();
 FILLCELL_X2 FILLER_22_1138 ();
 FILLCELL_X1 FILLER_22_1140 ();
 FILLCELL_X2 FILLER_22_1170 ();
 FILLCELL_X1 FILLER_22_1214 ();
 FILLCELL_X1 FILLER_22_1221 ();
 FILLCELL_X8 FILLER_22_1242 ();
 FILLCELL_X4 FILLER_22_1250 ();
 FILLCELL_X1 FILLER_22_1254 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X1 FILLER_23_402 ();
 FILLCELL_X2 FILLER_23_417 ();
 FILLCELL_X2 FILLER_23_426 ();
 FILLCELL_X1 FILLER_23_428 ();
 FILLCELL_X2 FILLER_23_436 ();
 FILLCELL_X1 FILLER_23_438 ();
 FILLCELL_X4 FILLER_23_456 ();
 FILLCELL_X1 FILLER_23_460 ();
 FILLCELL_X2 FILLER_23_470 ();
 FILLCELL_X4 FILLER_23_479 ();
 FILLCELL_X1 FILLER_23_483 ();
 FILLCELL_X2 FILLER_23_520 ();
 FILLCELL_X1 FILLER_23_522 ();
 FILLCELL_X4 FILLER_23_548 ();
 FILLCELL_X1 FILLER_23_552 ();
 FILLCELL_X2 FILLER_23_568 ();
 FILLCELL_X2 FILLER_23_576 ();
 FILLCELL_X1 FILLER_23_581 ();
 FILLCELL_X8 FILLER_23_593 ();
 FILLCELL_X4 FILLER_23_601 ();
 FILLCELL_X1 FILLER_23_605 ();
 FILLCELL_X4 FILLER_23_610 ();
 FILLCELL_X1 FILLER_23_626 ();
 FILLCELL_X8 FILLER_23_636 ();
 FILLCELL_X4 FILLER_23_644 ();
 FILLCELL_X2 FILLER_23_648 ();
 FILLCELL_X1 FILLER_23_650 ();
 FILLCELL_X8 FILLER_23_671 ();
 FILLCELL_X4 FILLER_23_708 ();
 FILLCELL_X2 FILLER_23_712 ();
 FILLCELL_X1 FILLER_23_721 ();
 FILLCELL_X4 FILLER_23_740 ();
 FILLCELL_X1 FILLER_23_744 ();
 FILLCELL_X1 FILLER_23_752 ();
 FILLCELL_X1 FILLER_23_757 ();
 FILLCELL_X1 FILLER_23_762 ();
 FILLCELL_X1 FILLER_23_771 ();
 FILLCELL_X8 FILLER_23_774 ();
 FILLCELL_X4 FILLER_23_782 ();
 FILLCELL_X1 FILLER_23_786 ();
 FILLCELL_X4 FILLER_23_833 ();
 FILLCELL_X2 FILLER_23_837 ();
 FILLCELL_X1 FILLER_23_839 ();
 FILLCELL_X2 FILLER_23_847 ();
 FILLCELL_X1 FILLER_23_849 ();
 FILLCELL_X4 FILLER_23_886 ();
 FILLCELL_X2 FILLER_23_890 ();
 FILLCELL_X8 FILLER_23_908 ();
 FILLCELL_X2 FILLER_23_935 ();
 FILLCELL_X1 FILLER_23_959 ();
 FILLCELL_X1 FILLER_23_984 ();
 FILLCELL_X4 FILLER_23_990 ();
 FILLCELL_X1 FILLER_23_994 ();
 FILLCELL_X8 FILLER_23_1005 ();
 FILLCELL_X2 FILLER_23_1013 ();
 FILLCELL_X1 FILLER_23_1015 ();
 FILLCELL_X8 FILLER_23_1021 ();
 FILLCELL_X4 FILLER_23_1029 ();
 FILLCELL_X1 FILLER_23_1033 ();
 FILLCELL_X2 FILLER_23_1041 ();
 FILLCELL_X2 FILLER_23_1050 ();
 FILLCELL_X1 FILLER_23_1052 ();
 FILLCELL_X16 FILLER_23_1075 ();
 FILLCELL_X4 FILLER_23_1091 ();
 FILLCELL_X2 FILLER_23_1095 ();
 FILLCELL_X1 FILLER_23_1097 ();
 FILLCELL_X16 FILLER_23_1105 ();
 FILLCELL_X8 FILLER_23_1121 ();
 FILLCELL_X2 FILLER_23_1129 ();
 FILLCELL_X8 FILLER_23_1138 ();
 FILLCELL_X32 FILLER_23_1166 ();
 FILLCELL_X1 FILLER_23_1198 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X8 FILLER_24_385 ();
 FILLCELL_X4 FILLER_24_393 ();
 FILLCELL_X2 FILLER_24_414 ();
 FILLCELL_X1 FILLER_24_416 ();
 FILLCELL_X1 FILLER_24_434 ();
 FILLCELL_X16 FILLER_24_442 ();
 FILLCELL_X2 FILLER_24_458 ();
 FILLCELL_X1 FILLER_24_460 ();
 FILLCELL_X16 FILLER_24_468 ();
 FILLCELL_X1 FILLER_24_504 ();
 FILLCELL_X8 FILLER_24_519 ();
 FILLCELL_X4 FILLER_24_527 ();
 FILLCELL_X1 FILLER_24_531 ();
 FILLCELL_X8 FILLER_24_552 ();
 FILLCELL_X2 FILLER_24_565 ();
 FILLCELL_X2 FILLER_24_595 ();
 FILLCELL_X2 FILLER_24_600 ();
 FILLCELL_X1 FILLER_24_602 ();
 FILLCELL_X2 FILLER_24_623 ();
 FILLCELL_X1 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X16 FILLER_24_640 ();
 FILLCELL_X2 FILLER_24_670 ();
 FILLCELL_X1 FILLER_24_672 ();
 FILLCELL_X4 FILLER_24_676 ();
 FILLCELL_X2 FILLER_24_680 ();
 FILLCELL_X4 FILLER_24_704 ();
 FILLCELL_X1 FILLER_24_708 ();
 FILLCELL_X8 FILLER_24_715 ();
 FILLCELL_X4 FILLER_24_728 ();
 FILLCELL_X2 FILLER_24_732 ();
 FILLCELL_X1 FILLER_24_734 ();
 FILLCELL_X4 FILLER_24_738 ();
 FILLCELL_X2 FILLER_24_742 ();
 FILLCELL_X2 FILLER_24_748 ();
 FILLCELL_X8 FILLER_24_774 ();
 FILLCELL_X1 FILLER_24_782 ();
 FILLCELL_X4 FILLER_24_803 ();
 FILLCELL_X2 FILLER_24_807 ();
 FILLCELL_X8 FILLER_24_811 ();
 FILLCELL_X4 FILLER_24_819 ();
 FILLCELL_X1 FILLER_24_823 ();
 FILLCELL_X4 FILLER_24_851 ();
 FILLCELL_X2 FILLER_24_855 ();
 FILLCELL_X16 FILLER_24_868 ();
 FILLCELL_X2 FILLER_24_884 ();
 FILLCELL_X1 FILLER_24_886 ();
 FILLCELL_X2 FILLER_24_898 ();
 FILLCELL_X1 FILLER_24_922 ();
 FILLCELL_X4 FILLER_24_955 ();
 FILLCELL_X1 FILLER_24_959 ();
 FILLCELL_X1 FILLER_24_966 ();
 FILLCELL_X4 FILLER_24_994 ();
 FILLCELL_X1 FILLER_24_998 ();
 FILLCELL_X2 FILLER_24_1093 ();
 FILLCELL_X4 FILLER_24_1115 ();
 FILLCELL_X4 FILLER_24_1139 ();
 FILLCELL_X16 FILLER_24_1150 ();
 FILLCELL_X8 FILLER_24_1166 ();
 FILLCELL_X2 FILLER_24_1223 ();
 FILLCELL_X1 FILLER_24_1225 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X1 FILLER_25_417 ();
 FILLCELL_X8 FILLER_25_425 ();
 FILLCELL_X4 FILLER_25_433 ();
 FILLCELL_X2 FILLER_25_437 ();
 FILLCELL_X4 FILLER_25_456 ();
 FILLCELL_X1 FILLER_25_460 ();
 FILLCELL_X8 FILLER_25_478 ();
 FILLCELL_X2 FILLER_25_486 ();
 FILLCELL_X1 FILLER_25_488 ();
 FILLCELL_X4 FILLER_25_507 ();
 FILLCELL_X2 FILLER_25_511 ();
 FILLCELL_X1 FILLER_25_513 ();
 FILLCELL_X8 FILLER_25_522 ();
 FILLCELL_X2 FILLER_25_530 ();
 FILLCELL_X2 FILLER_25_562 ();
 FILLCELL_X1 FILLER_25_567 ();
 FILLCELL_X1 FILLER_25_571 ();
 FILLCELL_X1 FILLER_25_576 ();
 FILLCELL_X2 FILLER_25_585 ();
 FILLCELL_X2 FILLER_25_591 ();
 FILLCELL_X2 FILLER_25_600 ();
 FILLCELL_X1 FILLER_25_611 ();
 FILLCELL_X2 FILLER_25_616 ();
 FILLCELL_X1 FILLER_25_622 ();
 FILLCELL_X16 FILLER_25_637 ();
 FILLCELL_X8 FILLER_25_653 ();
 FILLCELL_X4 FILLER_25_661 ();
 FILLCELL_X1 FILLER_25_665 ();
 FILLCELL_X16 FILLER_25_684 ();
 FILLCELL_X1 FILLER_25_703 ();
 FILLCELL_X2 FILLER_25_726 ();
 FILLCELL_X2 FILLER_25_748 ();
 FILLCELL_X1 FILLER_25_750 ();
 FILLCELL_X2 FILLER_25_771 ();
 FILLCELL_X1 FILLER_25_773 ();
 FILLCELL_X1 FILLER_25_782 ();
 FILLCELL_X2 FILLER_25_796 ();
 FILLCELL_X1 FILLER_25_798 ();
 FILLCELL_X2 FILLER_25_805 ();
 FILLCELL_X16 FILLER_25_819 ();
 FILLCELL_X2 FILLER_25_835 ();
 FILLCELL_X8 FILLER_25_849 ();
 FILLCELL_X1 FILLER_25_857 ();
 FILLCELL_X4 FILLER_25_871 ();
 FILLCELL_X4 FILLER_25_896 ();
 FILLCELL_X2 FILLER_25_900 ();
 FILLCELL_X1 FILLER_25_902 ();
 FILLCELL_X2 FILLER_25_914 ();
 FILLCELL_X4 FILLER_25_921 ();
 FILLCELL_X2 FILLER_25_925 ();
 FILLCELL_X1 FILLER_25_936 ();
 FILLCELL_X1 FILLER_25_955 ();
 FILLCELL_X16 FILLER_25_983 ();
 FILLCELL_X4 FILLER_25_999 ();
 FILLCELL_X32 FILLER_25_1010 ();
 FILLCELL_X16 FILLER_25_1042 ();
 FILLCELL_X8 FILLER_25_1058 ();
 FILLCELL_X2 FILLER_25_1066 ();
 FILLCELL_X1 FILLER_25_1068 ();
 FILLCELL_X4 FILLER_25_1073 ();
 FILLCELL_X2 FILLER_25_1077 ();
 FILLCELL_X2 FILLER_25_1086 ();
 FILLCELL_X1 FILLER_25_1088 ();
 FILLCELL_X16 FILLER_25_1101 ();
 FILLCELL_X1 FILLER_25_1117 ();
 FILLCELL_X1 FILLER_25_1125 ();
 FILLCELL_X1 FILLER_25_1153 ();
 FILLCELL_X8 FILLER_25_1181 ();
 FILLCELL_X2 FILLER_25_1189 ();
 FILLCELL_X16 FILLER_25_1196 ();
 FILLCELL_X4 FILLER_25_1212 ();
 FILLCELL_X1 FILLER_25_1216 ();
 FILLCELL_X16 FILLER_25_1223 ();
 FILLCELL_X8 FILLER_25_1239 ();
 FILLCELL_X1 FILLER_25_1247 ();
 FILLCELL_X2 FILLER_25_1253 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X16 FILLER_26_385 ();
 FILLCELL_X2 FILLER_26_401 ();
 FILLCELL_X1 FILLER_26_403 ();
 FILLCELL_X1 FILLER_26_421 ();
 FILLCELL_X4 FILLER_26_429 ();
 FILLCELL_X16 FILLER_26_440 ();
 FILLCELL_X4 FILLER_26_456 ();
 FILLCELL_X2 FILLER_26_460 ();
 FILLCELL_X16 FILLER_26_469 ();
 FILLCELL_X4 FILLER_26_485 ();
 FILLCELL_X2 FILLER_26_489 ();
 FILLCELL_X1 FILLER_26_491 ();
 FILLCELL_X1 FILLER_26_511 ();
 FILLCELL_X1 FILLER_26_516 ();
 FILLCELL_X1 FILLER_26_522 ();
 FILLCELL_X2 FILLER_26_527 ();
 FILLCELL_X1 FILLER_26_533 ();
 FILLCELL_X1 FILLER_26_539 ();
 FILLCELL_X1 FILLER_26_561 ();
 FILLCELL_X1 FILLER_26_567 ();
 FILLCELL_X1 FILLER_26_581 ();
 FILLCELL_X1 FILLER_26_587 ();
 FILLCELL_X1 FILLER_26_592 ();
 FILLCELL_X1 FILLER_26_597 ();
 FILLCELL_X2 FILLER_26_603 ();
 FILLCELL_X1 FILLER_26_608 ();
 FILLCELL_X2 FILLER_26_613 ();
 FILLCELL_X2 FILLER_26_619 ();
 FILLCELL_X2 FILLER_26_624 ();
 FILLCELL_X8 FILLER_26_632 ();
 FILLCELL_X4 FILLER_26_640 ();
 FILLCELL_X2 FILLER_26_644 ();
 FILLCELL_X1 FILLER_26_646 ();
 FILLCELL_X2 FILLER_26_672 ();
 FILLCELL_X2 FILLER_26_694 ();
 FILLCELL_X2 FILLER_26_700 ();
 FILLCELL_X16 FILLER_26_707 ();
 FILLCELL_X8 FILLER_26_723 ();
 FILLCELL_X4 FILLER_26_731 ();
 FILLCELL_X2 FILLER_26_757 ();
 FILLCELL_X1 FILLER_26_759 ();
 FILLCELL_X4 FILLER_26_763 ();
 FILLCELL_X1 FILLER_26_767 ();
 FILLCELL_X8 FILLER_26_773 ();
 FILLCELL_X1 FILLER_26_786 ();
 FILLCELL_X4 FILLER_26_791 ();
 FILLCELL_X2 FILLER_26_804 ();
 FILLCELL_X1 FILLER_26_806 ();
 FILLCELL_X2 FILLER_26_829 ();
 FILLCELL_X1 FILLER_26_831 ();
 FILLCELL_X2 FILLER_26_839 ();
 FILLCELL_X1 FILLER_26_841 ();
 FILLCELL_X8 FILLER_26_880 ();
 FILLCELL_X2 FILLER_26_888 ();
 FILLCELL_X2 FILLER_26_904 ();
 FILLCELL_X1 FILLER_26_906 ();
 FILLCELL_X4 FILLER_26_911 ();
 FILLCELL_X1 FILLER_26_915 ();
 FILLCELL_X2 FILLER_26_919 ();
 FILLCELL_X4 FILLER_26_928 ();
 FILLCELL_X8 FILLER_26_937 ();
 FILLCELL_X4 FILLER_26_945 ();
 FILLCELL_X2 FILLER_26_949 ();
 FILLCELL_X1 FILLER_26_951 ();
 FILLCELL_X8 FILLER_26_954 ();
 FILLCELL_X4 FILLER_26_962 ();
 FILLCELL_X1 FILLER_26_966 ();
 FILLCELL_X16 FILLER_26_977 ();
 FILLCELL_X4 FILLER_26_1022 ();
 FILLCELL_X2 FILLER_26_1026 ();
 FILLCELL_X1 FILLER_26_1034 ();
 FILLCELL_X1 FILLER_26_1040 ();
 FILLCELL_X2 FILLER_26_1047 ();
 FILLCELL_X2 FILLER_26_1054 ();
 FILLCELL_X2 FILLER_26_1076 ();
 FILLCELL_X1 FILLER_26_1078 ();
 FILLCELL_X16 FILLER_26_1099 ();
 FILLCELL_X4 FILLER_26_1115 ();
 FILLCELL_X4 FILLER_26_1133 ();
 FILLCELL_X1 FILLER_26_1137 ();
 FILLCELL_X16 FILLER_26_1152 ();
 FILLCELL_X1 FILLER_26_1184 ();
 FILLCELL_X2 FILLER_26_1190 ();
 FILLCELL_X2 FILLER_26_1195 ();
 FILLCELL_X1 FILLER_26_1197 ();
 FILLCELL_X1 FILLER_26_1205 ();
 FILLCELL_X1 FILLER_26_1221 ();
 FILLCELL_X1 FILLER_26_1227 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X16 FILLER_27_385 ();
 FILLCELL_X8 FILLER_27_401 ();
 FILLCELL_X4 FILLER_27_409 ();
 FILLCELL_X1 FILLER_27_413 ();
 FILLCELL_X8 FILLER_27_438 ();
 FILLCELL_X16 FILLER_27_467 ();
 FILLCELL_X8 FILLER_27_483 ();
 FILLCELL_X4 FILLER_27_491 ();
 FILLCELL_X2 FILLER_27_495 ();
 FILLCELL_X1 FILLER_27_506 ();
 FILLCELL_X1 FILLER_27_514 ();
 FILLCELL_X2 FILLER_27_526 ();
 FILLCELL_X2 FILLER_27_533 ();
 FILLCELL_X1 FILLER_27_539 ();
 FILLCELL_X16 FILLER_27_542 ();
 FILLCELL_X4 FILLER_27_558 ();
 FILLCELL_X2 FILLER_27_562 ();
 FILLCELL_X2 FILLER_27_591 ();
 FILLCELL_X2 FILLER_27_596 ();
 FILLCELL_X4 FILLER_27_602 ();
 FILLCELL_X1 FILLER_27_610 ();
 FILLCELL_X1 FILLER_27_618 ();
 FILLCELL_X16 FILLER_27_634 ();
 FILLCELL_X2 FILLER_27_650 ();
 FILLCELL_X2 FILLER_27_659 ();
 FILLCELL_X1 FILLER_27_677 ();
 FILLCELL_X16 FILLER_27_695 ();
 FILLCELL_X4 FILLER_27_711 ();
 FILLCELL_X2 FILLER_27_715 ();
 FILLCELL_X16 FILLER_27_743 ();
 FILLCELL_X1 FILLER_27_759 ();
 FILLCELL_X1 FILLER_27_776 ();
 FILLCELL_X1 FILLER_27_780 ();
 FILLCELL_X1 FILLER_27_785 ();
 FILLCELL_X1 FILLER_27_792 ();
 FILLCELL_X1 FILLER_27_797 ();
 FILLCELL_X2 FILLER_27_802 ();
 FILLCELL_X8 FILLER_27_817 ();
 FILLCELL_X4 FILLER_27_825 ();
 FILLCELL_X2 FILLER_27_829 ();
 FILLCELL_X1 FILLER_27_831 ();
 FILLCELL_X4 FILLER_27_841 ();
 FILLCELL_X2 FILLER_27_845 ();
 FILLCELL_X1 FILLER_27_847 ();
 FILLCELL_X4 FILLER_27_854 ();
 FILLCELL_X2 FILLER_27_858 ();
 FILLCELL_X4 FILLER_27_869 ();
 FILLCELL_X2 FILLER_27_873 ();
 FILLCELL_X2 FILLER_27_889 ();
 FILLCELL_X1 FILLER_27_891 ();
 FILLCELL_X1 FILLER_27_897 ();
 FILLCELL_X2 FILLER_27_901 ();
 FILLCELL_X1 FILLER_27_903 ();
 FILLCELL_X4 FILLER_27_911 ();
 FILLCELL_X2 FILLER_27_929 ();
 FILLCELL_X1 FILLER_27_934 ();
 FILLCELL_X4 FILLER_27_949 ();
 FILLCELL_X2 FILLER_27_953 ();
 FILLCELL_X4 FILLER_27_977 ();
 FILLCELL_X2 FILLER_27_981 ();
 FILLCELL_X1 FILLER_27_983 ();
 FILLCELL_X2 FILLER_27_989 ();
 FILLCELL_X2 FILLER_27_1012 ();
 FILLCELL_X2 FILLER_27_1041 ();
 FILLCELL_X1 FILLER_27_1043 ();
 FILLCELL_X1 FILLER_27_1062 ();
 FILLCELL_X4 FILLER_27_1074 ();
 FILLCELL_X2 FILLER_27_1078 ();
 FILLCELL_X1 FILLER_27_1080 ();
 FILLCELL_X8 FILLER_27_1086 ();
 FILLCELL_X1 FILLER_27_1094 ();
 FILLCELL_X8 FILLER_27_1117 ();
 FILLCELL_X2 FILLER_27_1125 ();
 FILLCELL_X1 FILLER_27_1134 ();
 FILLCELL_X2 FILLER_27_1169 ();
 FILLCELL_X2 FILLER_27_1180 ();
 FILLCELL_X4 FILLER_27_1189 ();
 FILLCELL_X2 FILLER_27_1193 ();
 FILLCELL_X4 FILLER_27_1202 ();
 FILLCELL_X2 FILLER_27_1206 ();
 FILLCELL_X4 FILLER_27_1222 ();
 FILLCELL_X2 FILLER_27_1226 ();
 FILLCELL_X1 FILLER_27_1228 ();
 FILLCELL_X1 FILLER_27_1247 ();
 FILLCELL_X4 FILLER_27_1251 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X16 FILLER_28_417 ();
 FILLCELL_X8 FILLER_28_433 ();
 FILLCELL_X2 FILLER_28_441 ();
 FILLCELL_X1 FILLER_28_443 ();
 FILLCELL_X16 FILLER_28_478 ();
 FILLCELL_X2 FILLER_28_494 ();
 FILLCELL_X1 FILLER_28_496 ();
 FILLCELL_X1 FILLER_28_527 ();
 FILLCELL_X1 FILLER_28_548 ();
 FILLCELL_X8 FILLER_28_572 ();
 FILLCELL_X2 FILLER_28_580 ();
 FILLCELL_X1 FILLER_28_582 ();
 FILLCELL_X1 FILLER_28_600 ();
 FILLCELL_X1 FILLER_28_606 ();
 FILLCELL_X1 FILLER_28_611 ();
 FILLCELL_X1 FILLER_28_618 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X1 FILLER_28_632 ();
 FILLCELL_X8 FILLER_28_674 ();
 FILLCELL_X8 FILLER_28_701 ();
 FILLCELL_X4 FILLER_28_709 ();
 FILLCELL_X2 FILLER_28_773 ();
 FILLCELL_X1 FILLER_28_775 ();
 FILLCELL_X8 FILLER_28_794 ();
 FILLCELL_X2 FILLER_28_802 ();
 FILLCELL_X2 FILLER_28_857 ();
 FILLCELL_X1 FILLER_28_863 ();
 FILLCELL_X4 FILLER_28_884 ();
 FILLCELL_X2 FILLER_28_888 ();
 FILLCELL_X2 FILLER_28_892 ();
 FILLCELL_X2 FILLER_28_908 ();
 FILLCELL_X1 FILLER_28_910 ();
 FILLCELL_X1 FILLER_28_914 ();
 FILLCELL_X2 FILLER_28_920 ();
 FILLCELL_X1 FILLER_28_922 ();
 FILLCELL_X8 FILLER_28_930 ();
 FILLCELL_X2 FILLER_28_938 ();
 FILLCELL_X8 FILLER_28_947 ();
 FILLCELL_X16 FILLER_28_962 ();
 FILLCELL_X4 FILLER_28_978 ();
 FILLCELL_X1 FILLER_28_982 ();
 FILLCELL_X2 FILLER_28_1010 ();
 FILLCELL_X1 FILLER_28_1012 ();
 FILLCELL_X8 FILLER_28_1020 ();
 FILLCELL_X4 FILLER_28_1028 ();
 FILLCELL_X1 FILLER_28_1032 ();
 FILLCELL_X4 FILLER_28_1060 ();
 FILLCELL_X1 FILLER_28_1064 ();
 FILLCELL_X2 FILLER_28_1087 ();
 FILLCELL_X1 FILLER_28_1089 ();
 FILLCELL_X4 FILLER_28_1117 ();
 FILLCELL_X2 FILLER_28_1121 ();
 FILLCELL_X1 FILLER_28_1123 ();
 FILLCELL_X2 FILLER_28_1140 ();
 FILLCELL_X1 FILLER_28_1142 ();
 FILLCELL_X4 FILLER_28_1150 ();
 FILLCELL_X1 FILLER_28_1154 ();
 FILLCELL_X1 FILLER_28_1191 ();
 FILLCELL_X32 FILLER_28_1197 ();
 FILLCELL_X2 FILLER_28_1229 ();
 FILLCELL_X8 FILLER_28_1247 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X16 FILLER_29_449 ();
 FILLCELL_X4 FILLER_29_465 ();
 FILLCELL_X1 FILLER_29_469 ();
 FILLCELL_X16 FILLER_29_478 ();
 FILLCELL_X2 FILLER_29_514 ();
 FILLCELL_X1 FILLER_29_516 ();
 FILLCELL_X4 FILLER_29_521 ();
 FILLCELL_X2 FILLER_29_525 ();
 FILLCELL_X1 FILLER_29_527 ();
 FILLCELL_X2 FILLER_29_546 ();
 FILLCELL_X1 FILLER_29_548 ();
 FILLCELL_X2 FILLER_29_582 ();
 FILLCELL_X1 FILLER_29_588 ();
 FILLCELL_X4 FILLER_29_592 ();
 FILLCELL_X1 FILLER_29_602 ();
 FILLCELL_X1 FILLER_29_607 ();
 FILLCELL_X2 FILLER_29_620 ();
 FILLCELL_X1 FILLER_29_622 ();
 FILLCELL_X2 FILLER_29_627 ();
 FILLCELL_X2 FILLER_29_640 ();
 FILLCELL_X1 FILLER_29_642 ();
 FILLCELL_X8 FILLER_29_650 ();
 FILLCELL_X2 FILLER_29_658 ();
 FILLCELL_X1 FILLER_29_660 ();
 FILLCELL_X4 FILLER_29_685 ();
 FILLCELL_X1 FILLER_29_689 ();
 FILLCELL_X8 FILLER_29_694 ();
 FILLCELL_X4 FILLER_29_702 ();
 FILLCELL_X2 FILLER_29_706 ();
 FILLCELL_X8 FILLER_29_715 ();
 FILLCELL_X4 FILLER_29_723 ();
 FILLCELL_X1 FILLER_29_727 ();
 FILLCELL_X8 FILLER_29_737 ();
 FILLCELL_X4 FILLER_29_745 ();
 FILLCELL_X1 FILLER_29_749 ();
 FILLCELL_X1 FILLER_29_772 ();
 FILLCELL_X2 FILLER_29_777 ();
 FILLCELL_X1 FILLER_29_799 ();
 FILLCELL_X2 FILLER_29_803 ();
 FILLCELL_X8 FILLER_29_823 ();
 FILLCELL_X1 FILLER_29_831 ();
 FILLCELL_X2 FILLER_29_864 ();
 FILLCELL_X1 FILLER_29_866 ();
 FILLCELL_X8 FILLER_29_873 ();
 FILLCELL_X2 FILLER_29_881 ();
 FILLCELL_X1 FILLER_29_883 ();
 FILLCELL_X2 FILLER_29_889 ();
 FILLCELL_X1 FILLER_29_891 ();
 FILLCELL_X2 FILLER_29_895 ();
 FILLCELL_X1 FILLER_29_897 ();
 FILLCELL_X1 FILLER_29_912 ();
 FILLCELL_X4 FILLER_29_961 ();
 FILLCELL_X8 FILLER_29_992 ();
 FILLCELL_X2 FILLER_29_1000 ();
 FILLCELL_X4 FILLER_29_1007 ();
 FILLCELL_X1 FILLER_29_1011 ();
 FILLCELL_X8 FILLER_29_1020 ();
 FILLCELL_X1 FILLER_29_1028 ();
 FILLCELL_X4 FILLER_29_1039 ();
 FILLCELL_X2 FILLER_29_1043 ();
 FILLCELL_X1 FILLER_29_1045 ();
 FILLCELL_X2 FILLER_29_1050 ();
 FILLCELL_X1 FILLER_29_1052 ();
 FILLCELL_X4 FILLER_29_1056 ();
 FILLCELL_X2 FILLER_29_1060 ();
 FILLCELL_X1 FILLER_29_1062 ();
 FILLCELL_X8 FILLER_29_1070 ();
 FILLCELL_X1 FILLER_29_1090 ();
 FILLCELL_X4 FILLER_29_1097 ();
 FILLCELL_X2 FILLER_29_1101 ();
 FILLCELL_X8 FILLER_29_1112 ();
 FILLCELL_X4 FILLER_29_1120 ();
 FILLCELL_X2 FILLER_29_1124 ();
 FILLCELL_X1 FILLER_29_1126 ();
 FILLCELL_X4 FILLER_29_1132 ();
 FILLCELL_X1 FILLER_29_1136 ();
 FILLCELL_X2 FILLER_29_1157 ();
 FILLCELL_X1 FILLER_29_1159 ();
 FILLCELL_X1 FILLER_29_1174 ();
 FILLCELL_X1 FILLER_29_1182 ();
 FILLCELL_X2 FILLER_29_1203 ();
 FILLCELL_X2 FILLER_29_1232 ();
 FILLCELL_X1 FILLER_29_1234 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X16 FILLER_30_225 ();
 FILLCELL_X8 FILLER_30_241 ();
 FILLCELL_X4 FILLER_30_249 ();
 FILLCELL_X1 FILLER_30_253 ();
 FILLCELL_X16 FILLER_30_257 ();
 FILLCELL_X1 FILLER_30_293 ();
 FILLCELL_X16 FILLER_30_301 ();
 FILLCELL_X1 FILLER_30_321 ();
 FILLCELL_X4 FILLER_30_325 ();
 FILLCELL_X1 FILLER_30_329 ();
 FILLCELL_X4 FILLER_30_334 ();
 FILLCELL_X2 FILLER_30_338 ();
 FILLCELL_X2 FILLER_30_343 ();
 FILLCELL_X1 FILLER_30_345 ();
 FILLCELL_X8 FILLER_30_367 ();
 FILLCELL_X4 FILLER_30_375 ();
 FILLCELL_X8 FILLER_30_383 ();
 FILLCELL_X1 FILLER_30_391 ();
 FILLCELL_X8 FILLER_30_419 ();
 FILLCELL_X32 FILLER_30_434 ();
 FILLCELL_X4 FILLER_30_466 ();
 FILLCELL_X1 FILLER_30_470 ();
 FILLCELL_X8 FILLER_30_491 ();
 FILLCELL_X2 FILLER_30_499 ();
 FILLCELL_X1 FILLER_30_501 ();
 FILLCELL_X1 FILLER_30_524 ();
 FILLCELL_X1 FILLER_30_529 ();
 FILLCELL_X1 FILLER_30_544 ();
 FILLCELL_X1 FILLER_30_554 ();
 FILLCELL_X2 FILLER_30_558 ();
 FILLCELL_X2 FILLER_30_575 ();
 FILLCELL_X4 FILLER_30_580 ();
 FILLCELL_X2 FILLER_30_584 ();
 FILLCELL_X1 FILLER_30_593 ();
 FILLCELL_X1 FILLER_30_608 ();
 FILLCELL_X4 FILLER_30_616 ();
 FILLCELL_X1 FILLER_30_620 ();
 FILLCELL_X4 FILLER_30_624 ();
 FILLCELL_X2 FILLER_30_628 ();
 FILLCELL_X1 FILLER_30_630 ();
 FILLCELL_X1 FILLER_30_632 ();
 FILLCELL_X8 FILLER_30_637 ();
 FILLCELL_X16 FILLER_30_662 ();
 FILLCELL_X8 FILLER_30_678 ();
 FILLCELL_X4 FILLER_30_686 ();
 FILLCELL_X8 FILLER_30_717 ();
 FILLCELL_X4 FILLER_30_725 ();
 FILLCELL_X1 FILLER_30_729 ();
 FILLCELL_X1 FILLER_30_771 ();
 FILLCELL_X1 FILLER_30_776 ();
 FILLCELL_X1 FILLER_30_781 ();
 FILLCELL_X2 FILLER_30_786 ();
 FILLCELL_X2 FILLER_30_792 ();
 FILLCELL_X2 FILLER_30_803 ();
 FILLCELL_X4 FILLER_30_823 ();
 FILLCELL_X1 FILLER_30_827 ();
 FILLCELL_X4 FILLER_30_834 ();
 FILLCELL_X1 FILLER_30_842 ();
 FILLCELL_X2 FILLER_30_854 ();
 FILLCELL_X2 FILLER_30_864 ();
 FILLCELL_X4 FILLER_30_886 ();
 FILLCELL_X2 FILLER_30_906 ();
 FILLCELL_X1 FILLER_30_908 ();
 FILLCELL_X2 FILLER_30_930 ();
 FILLCELL_X4 FILLER_30_972 ();
 FILLCELL_X2 FILLER_30_976 ();
 FILLCELL_X4 FILLER_30_1009 ();
 FILLCELL_X2 FILLER_30_1013 ();
 FILLCELL_X2 FILLER_30_1076 ();
 FILLCELL_X1 FILLER_30_1078 ();
 FILLCELL_X2 FILLER_30_1099 ();
 FILLCELL_X16 FILLER_30_1142 ();
 FILLCELL_X4 FILLER_30_1158 ();
 FILLCELL_X2 FILLER_30_1169 ();
 FILLCELL_X1 FILLER_30_1223 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X8 FILLER_31_225 ();
 FILLCELL_X2 FILLER_31_233 ();
 FILLCELL_X2 FILLER_31_242 ();
 FILLCELL_X1 FILLER_31_244 ();
 FILLCELL_X4 FILLER_31_278 ();
 FILLCELL_X2 FILLER_31_345 ();
 FILLCELL_X2 FILLER_31_380 ();
 FILLCELL_X1 FILLER_31_382 ();
 FILLCELL_X4 FILLER_31_410 ();
 FILLCELL_X2 FILLER_31_414 ();
 FILLCELL_X8 FILLER_31_419 ();
 FILLCELL_X4 FILLER_31_427 ();
 FILLCELL_X16 FILLER_31_451 ();
 FILLCELL_X1 FILLER_31_467 ();
 FILLCELL_X4 FILLER_31_475 ();
 FILLCELL_X1 FILLER_31_479 ();
 FILLCELL_X2 FILLER_31_521 ();
 FILLCELL_X2 FILLER_31_532 ();
 FILLCELL_X1 FILLER_31_534 ();
 FILLCELL_X1 FILLER_31_557 ();
 FILLCELL_X2 FILLER_31_561 ();
 FILLCELL_X8 FILLER_31_567 ();
 FILLCELL_X1 FILLER_31_575 ();
 FILLCELL_X1 FILLER_31_583 ();
 FILLCELL_X2 FILLER_31_616 ();
 FILLCELL_X32 FILLER_31_630 ();
 FILLCELL_X4 FILLER_31_662 ();
 FILLCELL_X4 FILLER_31_671 ();
 FILLCELL_X32 FILLER_31_682 ();
 FILLCELL_X8 FILLER_31_714 ();
 FILLCELL_X1 FILLER_31_722 ();
 FILLCELL_X2 FILLER_31_743 ();
 FILLCELL_X1 FILLER_31_745 ();
 FILLCELL_X4 FILLER_31_763 ();
 FILLCELL_X2 FILLER_31_797 ();
 FILLCELL_X1 FILLER_31_799 ();
 FILLCELL_X2 FILLER_31_806 ();
 FILLCELL_X1 FILLER_31_808 ();
 FILLCELL_X4 FILLER_31_822 ();
 FILLCELL_X2 FILLER_31_826 ();
 FILLCELL_X8 FILLER_31_836 ();
 FILLCELL_X1 FILLER_31_844 ();
 FILLCELL_X16 FILLER_31_859 ();
 FILLCELL_X8 FILLER_31_878 ();
 FILLCELL_X4 FILLER_31_886 ();
 FILLCELL_X2 FILLER_31_890 ();
 FILLCELL_X2 FILLER_31_903 ();
 FILLCELL_X1 FILLER_31_905 ();
 FILLCELL_X2 FILLER_31_909 ();
 FILLCELL_X16 FILLER_31_933 ();
 FILLCELL_X8 FILLER_31_949 ();
 FILLCELL_X4 FILLER_31_957 ();
 FILLCELL_X2 FILLER_31_961 ();
 FILLCELL_X1 FILLER_31_963 ();
 FILLCELL_X8 FILLER_31_986 ();
 FILLCELL_X2 FILLER_31_994 ();
 FILLCELL_X4 FILLER_31_1027 ();
 FILLCELL_X2 FILLER_31_1031 ();
 FILLCELL_X16 FILLER_31_1038 ();
 FILLCELL_X8 FILLER_31_1054 ();
 FILLCELL_X4 FILLER_31_1067 ();
 FILLCELL_X1 FILLER_31_1071 ();
 FILLCELL_X16 FILLER_31_1086 ();
 FILLCELL_X16 FILLER_31_1115 ();
 FILLCELL_X8 FILLER_31_1131 ();
 FILLCELL_X1 FILLER_31_1139 ();
 FILLCELL_X4 FILLER_31_1156 ();
 FILLCELL_X2 FILLER_31_1177 ();
 FILLCELL_X1 FILLER_31_1189 ();
 FILLCELL_X8 FILLER_31_1195 ();
 FILLCELL_X2 FILLER_31_1203 ();
 FILLCELL_X1 FILLER_31_1205 ();
 FILLCELL_X8 FILLER_31_1213 ();
 FILLCELL_X2 FILLER_31_1221 ();
 FILLCELL_X1 FILLER_31_1227 ();
 FILLCELL_X2 FILLER_31_1235 ();
 FILLCELL_X2 FILLER_31_1244 ();
 FILLCELL_X2 FILLER_31_1252 ();
 FILLCELL_X1 FILLER_31_1254 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X16 FILLER_32_193 ();
 FILLCELL_X8 FILLER_32_209 ();
 FILLCELL_X1 FILLER_32_217 ();
 FILLCELL_X8 FILLER_32_262 ();
 FILLCELL_X4 FILLER_32_315 ();
 FILLCELL_X1 FILLER_32_323 ();
 FILLCELL_X8 FILLER_32_327 ();
 FILLCELL_X4 FILLER_32_340 ();
 FILLCELL_X2 FILLER_32_349 ();
 FILLCELL_X1 FILLER_32_351 ();
 FILLCELL_X4 FILLER_32_395 ();
 FILLCELL_X1 FILLER_32_411 ();
 FILLCELL_X1 FILLER_32_416 ();
 FILLCELL_X4 FILLER_32_437 ();
 FILLCELL_X2 FILLER_32_441 ();
 FILLCELL_X16 FILLER_32_450 ();
 FILLCELL_X4 FILLER_32_466 ();
 FILLCELL_X1 FILLER_32_470 ();
 FILLCELL_X8 FILLER_32_478 ();
 FILLCELL_X1 FILLER_32_506 ();
 FILLCELL_X8 FILLER_32_534 ();
 FILLCELL_X4 FILLER_32_542 ();
 FILLCELL_X2 FILLER_32_546 ();
 FILLCELL_X1 FILLER_32_548 ();
 FILLCELL_X1 FILLER_32_561 ();
 FILLCELL_X2 FILLER_32_566 ();
 FILLCELL_X4 FILLER_32_575 ();
 FILLCELL_X1 FILLER_32_579 ();
 FILLCELL_X4 FILLER_32_594 ();
 FILLCELL_X1 FILLER_32_598 ();
 FILLCELL_X2 FILLER_32_607 ();
 FILLCELL_X1 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_617 ();
 FILLCELL_X2 FILLER_32_621 ();
 FILLCELL_X1 FILLER_32_623 ();
 FILLCELL_X1 FILLER_32_649 ();
 FILLCELL_X16 FILLER_32_704 ();
 FILLCELL_X4 FILLER_32_720 ();
 FILLCELL_X4 FILLER_32_753 ();
 FILLCELL_X1 FILLER_32_757 ();
 FILLCELL_X2 FILLER_32_767 ();
 FILLCELL_X2 FILLER_32_772 ();
 FILLCELL_X2 FILLER_32_776 ();
 FILLCELL_X1 FILLER_32_778 ();
 FILLCELL_X1 FILLER_32_784 ();
 FILLCELL_X2 FILLER_32_790 ();
 FILLCELL_X1 FILLER_32_801 ();
 FILLCELL_X4 FILLER_32_810 ();
 FILLCELL_X1 FILLER_32_814 ();
 FILLCELL_X4 FILLER_32_835 ();
 FILLCELL_X1 FILLER_32_841 ();
 FILLCELL_X2 FILLER_32_844 ();
 FILLCELL_X4 FILLER_32_866 ();
 FILLCELL_X2 FILLER_32_870 ();
 FILLCELL_X1 FILLER_32_872 ();
 FILLCELL_X8 FILLER_32_894 ();
 FILLCELL_X1 FILLER_32_902 ();
 FILLCELL_X1 FILLER_32_919 ();
 FILLCELL_X4 FILLER_32_927 ();
 FILLCELL_X2 FILLER_32_931 ();
 FILLCELL_X1 FILLER_32_933 ();
 FILLCELL_X1 FILLER_32_954 ();
 FILLCELL_X1 FILLER_32_962 ();
 FILLCELL_X4 FILLER_32_975 ();
 FILLCELL_X2 FILLER_32_994 ();
 FILLCELL_X16 FILLER_32_1003 ();
 FILLCELL_X4 FILLER_32_1026 ();
 FILLCELL_X2 FILLER_32_1030 ();
 FILLCELL_X1 FILLER_32_1032 ();
 FILLCELL_X8 FILLER_32_1082 ();
 FILLCELL_X1 FILLER_32_1090 ();
 FILLCELL_X8 FILLER_32_1104 ();
 FILLCELL_X4 FILLER_32_1112 ();
 FILLCELL_X2 FILLER_32_1116 ();
 FILLCELL_X1 FILLER_32_1118 ();
 FILLCELL_X1 FILLER_32_1168 ();
 FILLCELL_X1 FILLER_32_1178 ();
 FILLCELL_X1 FILLER_32_1186 ();
 FILLCELL_X1 FILLER_32_1207 ();
 FILLCELL_X4 FILLER_32_1213 ();
 FILLCELL_X2 FILLER_32_1217 ();
 FILLCELL_X1 FILLER_32_1219 ();
 FILLCELL_X2 FILLER_32_1233 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_161 ();
 FILLCELL_X4 FILLER_33_169 ();
 FILLCELL_X2 FILLER_33_173 ();
 FILLCELL_X8 FILLER_33_195 ();
 FILLCELL_X4 FILLER_33_203 ();
 FILLCELL_X2 FILLER_33_230 ();
 FILLCELL_X2 FILLER_33_236 ();
 FILLCELL_X8 FILLER_33_241 ();
 FILLCELL_X4 FILLER_33_249 ();
 FILLCELL_X2 FILLER_33_269 ();
 FILLCELL_X2 FILLER_33_331 ();
 FILLCELL_X2 FILLER_33_342 ();
 FILLCELL_X4 FILLER_33_347 ();
 FILLCELL_X1 FILLER_33_351 ();
 FILLCELL_X4 FILLER_33_381 ();
 FILLCELL_X2 FILLER_33_389 ();
 FILLCELL_X8 FILLER_33_414 ();
 FILLCELL_X4 FILLER_33_422 ();
 FILLCELL_X1 FILLER_33_426 ();
 FILLCELL_X2 FILLER_33_447 ();
 FILLCELL_X1 FILLER_33_474 ();
 FILLCELL_X8 FILLER_33_487 ();
 FILLCELL_X2 FILLER_33_495 ();
 FILLCELL_X1 FILLER_33_497 ();
 FILLCELL_X2 FILLER_33_523 ();
 FILLCELL_X1 FILLER_33_525 ();
 FILLCELL_X2 FILLER_33_551 ();
 FILLCELL_X1 FILLER_33_553 ();
 FILLCELL_X2 FILLER_33_588 ();
 FILLCELL_X1 FILLER_33_590 ();
 FILLCELL_X4 FILLER_33_605 ();
 FILLCELL_X1 FILLER_33_609 ();
 FILLCELL_X8 FILLER_33_627 ();
 FILLCELL_X4 FILLER_33_635 ();
 FILLCELL_X8 FILLER_33_670 ();
 FILLCELL_X2 FILLER_33_678 ();
 FILLCELL_X2 FILLER_33_690 ();
 FILLCELL_X1 FILLER_33_692 ();
 FILLCELL_X1 FILLER_33_725 ();
 FILLCELL_X8 FILLER_33_735 ();
 FILLCELL_X16 FILLER_33_747 ();
 FILLCELL_X2 FILLER_33_763 ();
 FILLCELL_X4 FILLER_33_772 ();
 FILLCELL_X2 FILLER_33_776 ();
 FILLCELL_X4 FILLER_33_788 ();
 FILLCELL_X2 FILLER_33_792 ();
 FILLCELL_X1 FILLER_33_798 ();
 FILLCELL_X8 FILLER_33_815 ();
 FILLCELL_X2 FILLER_33_823 ();
 FILLCELL_X2 FILLER_33_828 ();
 FILLCELL_X4 FILLER_33_835 ();
 FILLCELL_X2 FILLER_33_839 ();
 FILLCELL_X1 FILLER_33_841 ();
 FILLCELL_X16 FILLER_33_851 ();
 FILLCELL_X1 FILLER_33_867 ();
 FILLCELL_X2 FILLER_33_884 ();
 FILLCELL_X1 FILLER_33_886 ();
 FILLCELL_X2 FILLER_33_897 ();
 FILLCELL_X1 FILLER_33_899 ();
 FILLCELL_X1 FILLER_33_913 ();
 FILLCELL_X16 FILLER_33_921 ();
 FILLCELL_X8 FILLER_33_937 ();
 FILLCELL_X4 FILLER_33_945 ();
 FILLCELL_X1 FILLER_33_949 ();
 FILLCELL_X4 FILLER_33_970 ();
 FILLCELL_X8 FILLER_33_1058 ();
 FILLCELL_X2 FILLER_33_1066 ();
 FILLCELL_X16 FILLER_33_1071 ();
 FILLCELL_X2 FILLER_33_1087 ();
 FILLCELL_X1 FILLER_33_1096 ();
 FILLCELL_X4 FILLER_33_1134 ();
 FILLCELL_X2 FILLER_33_1159 ();
 FILLCELL_X1 FILLER_33_1161 ();
 FILLCELL_X2 FILLER_33_1169 ();
 FILLCELL_X1 FILLER_33_1171 ();
 FILLCELL_X4 FILLER_33_1177 ();
 FILLCELL_X2 FILLER_33_1181 ();
 FILLCELL_X1 FILLER_33_1183 ();
 FILLCELL_X8 FILLER_33_1189 ();
 FILLCELL_X4 FILLER_33_1197 ();
 FILLCELL_X2 FILLER_33_1201 ();
 FILLCELL_X2 FILLER_33_1228 ();
 FILLCELL_X2 FILLER_33_1244 ();
 FILLCELL_X2 FILLER_33_1249 ();
 FILLCELL_X1 FILLER_33_1251 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X16 FILLER_34_97 ();
 FILLCELL_X1 FILLER_34_113 ();
 FILLCELL_X8 FILLER_34_141 ();
 FILLCELL_X4 FILLER_34_149 ();
 FILLCELL_X1 FILLER_34_153 ();
 FILLCELL_X8 FILLER_34_161 ();
 FILLCELL_X1 FILLER_34_169 ();
 FILLCELL_X16 FILLER_34_204 ();
 FILLCELL_X2 FILLER_34_292 ();
 FILLCELL_X16 FILLER_34_297 ();
 FILLCELL_X8 FILLER_34_313 ();
 FILLCELL_X4 FILLER_34_321 ();
 FILLCELL_X2 FILLER_34_325 ();
 FILLCELL_X1 FILLER_34_327 ();
 FILLCELL_X4 FILLER_34_368 ();
 FILLCELL_X1 FILLER_34_375 ();
 FILLCELL_X1 FILLER_34_399 ();
 FILLCELL_X4 FILLER_34_404 ();
 FILLCELL_X4 FILLER_34_432 ();
 FILLCELL_X2 FILLER_34_436 ();
 FILLCELL_X1 FILLER_34_438 ();
 FILLCELL_X2 FILLER_34_453 ();
 FILLCELL_X2 FILLER_34_475 ();
 FILLCELL_X2 FILLER_34_487 ();
 FILLCELL_X4 FILLER_34_496 ();
 FILLCELL_X8 FILLER_34_505 ();
 FILLCELL_X2 FILLER_34_513 ();
 FILLCELL_X1 FILLER_34_515 ();
 FILLCELL_X4 FILLER_34_530 ();
 FILLCELL_X2 FILLER_34_534 ();
 FILLCELL_X1 FILLER_34_536 ();
 FILLCELL_X8 FILLER_34_560 ();
 FILLCELL_X1 FILLER_34_568 ();
 FILLCELL_X4 FILLER_34_576 ();
 FILLCELL_X2 FILLER_34_614 ();
 FILLCELL_X1 FILLER_34_616 ();
 FILLCELL_X1 FILLER_34_624 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X4 FILLER_34_632 ();
 FILLCELL_X2 FILLER_34_636 ();
 FILLCELL_X2 FILLER_34_645 ();
 FILLCELL_X4 FILLER_34_702 ();
 FILLCELL_X1 FILLER_34_706 ();
 FILLCELL_X4 FILLER_34_711 ();
 FILLCELL_X1 FILLER_34_715 ();
 FILLCELL_X4 FILLER_34_736 ();
 FILLCELL_X2 FILLER_34_746 ();
 FILLCELL_X2 FILLER_34_785 ();
 FILLCELL_X8 FILLER_34_826 ();
 FILLCELL_X4 FILLER_34_834 ();
 FILLCELL_X2 FILLER_34_838 ();
 FILLCELL_X4 FILLER_34_851 ();
 FILLCELL_X4 FILLER_34_867 ();
 FILLCELL_X1 FILLER_34_871 ();
 FILLCELL_X2 FILLER_34_887 ();
 FILLCELL_X1 FILLER_34_889 ();
 FILLCELL_X4 FILLER_34_906 ();
 FILLCELL_X1 FILLER_34_910 ();
 FILLCELL_X2 FILLER_34_915 ();
 FILLCELL_X1 FILLER_34_917 ();
 FILLCELL_X2 FILLER_34_955 ();
 FILLCELL_X1 FILLER_34_957 ();
 FILLCELL_X1 FILLER_34_965 ();
 FILLCELL_X32 FILLER_34_979 ();
 FILLCELL_X4 FILLER_34_1016 ();
 FILLCELL_X1 FILLER_34_1020 ();
 FILLCELL_X1 FILLER_34_1030 ();
 FILLCELL_X1 FILLER_34_1038 ();
 FILLCELL_X1 FILLER_34_1043 ();
 FILLCELL_X1 FILLER_34_1051 ();
 FILLCELL_X4 FILLER_34_1085 ();
 FILLCELL_X4 FILLER_34_1113 ();
 FILLCELL_X2 FILLER_34_1117 ();
 FILLCELL_X1 FILLER_34_1119 ();
 FILLCELL_X4 FILLER_34_1129 ();
 FILLCELL_X2 FILLER_34_1133 ();
 FILLCELL_X4 FILLER_34_1150 ();
 FILLCELL_X1 FILLER_34_1154 ();
 FILLCELL_X4 FILLER_34_1219 ();
 FILLCELL_X1 FILLER_34_1223 ();
 FILLCELL_X4 FILLER_34_1232 ();
 FILLCELL_X1 FILLER_34_1236 ();
 FILLCELL_X1 FILLER_34_1248 ();
 FILLCELL_X2 FILLER_34_1253 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X4 FILLER_35_129 ();
 FILLCELL_X1 FILLER_35_133 ();
 FILLCELL_X2 FILLER_35_181 ();
 FILLCELL_X4 FILLER_35_237 ();
 FILLCELL_X1 FILLER_35_241 ();
 FILLCELL_X2 FILLER_35_260 ();
 FILLCELL_X1 FILLER_35_262 ();
 FILLCELL_X4 FILLER_35_273 ();
 FILLCELL_X2 FILLER_35_281 ();
 FILLCELL_X2 FILLER_35_296 ();
 FILLCELL_X4 FILLER_35_302 ();
 FILLCELL_X4 FILLER_35_309 ();
 FILLCELL_X2 FILLER_35_313 ();
 FILLCELL_X2 FILLER_35_324 ();
 FILLCELL_X4 FILLER_35_329 ();
 FILLCELL_X1 FILLER_35_333 ();
 FILLCELL_X8 FILLER_35_339 ();
 FILLCELL_X4 FILLER_35_347 ();
 FILLCELL_X2 FILLER_35_351 ();
 FILLCELL_X1 FILLER_35_353 ();
 FILLCELL_X4 FILLER_35_357 ();
 FILLCELL_X2 FILLER_35_361 ();
 FILLCELL_X8 FILLER_35_383 ();
 FILLCELL_X4 FILLER_35_391 ();
 FILLCELL_X1 FILLER_35_395 ();
 FILLCELL_X16 FILLER_35_416 ();
 FILLCELL_X2 FILLER_35_432 ();
 FILLCELL_X4 FILLER_35_441 ();
 FILLCELL_X2 FILLER_35_445 ();
 FILLCELL_X4 FILLER_35_465 ();
 FILLCELL_X1 FILLER_35_473 ();
 FILLCELL_X8 FILLER_35_500 ();
 FILLCELL_X1 FILLER_35_508 ();
 FILLCELL_X2 FILLER_35_525 ();
 FILLCELL_X1 FILLER_35_527 ();
 FILLCELL_X8 FILLER_35_535 ();
 FILLCELL_X8 FILLER_35_592 ();
 FILLCELL_X2 FILLER_35_600 ();
 FILLCELL_X1 FILLER_35_602 ();
 FILLCELL_X4 FILLER_35_610 ();
 FILLCELL_X2 FILLER_35_614 ();
 FILLCELL_X1 FILLER_35_616 ();
 FILLCELL_X2 FILLER_35_636 ();
 FILLCELL_X1 FILLER_35_655 ();
 FILLCELL_X16 FILLER_35_663 ();
 FILLCELL_X4 FILLER_35_679 ();
 FILLCELL_X2 FILLER_35_683 ();
 FILLCELL_X1 FILLER_35_685 ();
 FILLCELL_X4 FILLER_35_699 ();
 FILLCELL_X2 FILLER_35_703 ();
 FILLCELL_X1 FILLER_35_705 ();
 FILLCELL_X1 FILLER_35_725 ();
 FILLCELL_X4 FILLER_35_731 ();
 FILLCELL_X2 FILLER_35_735 ();
 FILLCELL_X2 FILLER_35_739 ();
 FILLCELL_X16 FILLER_35_752 ();
 FILLCELL_X8 FILLER_35_790 ();
 FILLCELL_X4 FILLER_35_798 ();
 FILLCELL_X8 FILLER_35_806 ();
 FILLCELL_X4 FILLER_35_814 ();
 FILLCELL_X1 FILLER_35_818 ();
 FILLCELL_X1 FILLER_35_828 ();
 FILLCELL_X16 FILLER_35_845 ();
 FILLCELL_X8 FILLER_35_861 ();
 FILLCELL_X2 FILLER_35_869 ();
 FILLCELL_X4 FILLER_35_878 ();
 FILLCELL_X2 FILLER_35_904 ();
 FILLCELL_X4 FILLER_35_923 ();
 FILLCELL_X1 FILLER_35_927 ();
 FILLCELL_X8 FILLER_35_933 ();
 FILLCELL_X2 FILLER_35_941 ();
 FILLCELL_X1 FILLER_35_943 ();
 FILLCELL_X4 FILLER_35_955 ();
 FILLCELL_X2 FILLER_35_959 ();
 FILLCELL_X1 FILLER_35_961 ();
 FILLCELL_X8 FILLER_35_974 ();
 FILLCELL_X2 FILLER_35_982 ();
 FILLCELL_X1 FILLER_35_984 ();
 FILLCELL_X4 FILLER_35_1005 ();
 FILLCELL_X2 FILLER_35_1009 ();
 FILLCELL_X1 FILLER_35_1011 ();
 FILLCELL_X2 FILLER_35_1023 ();
 FILLCELL_X4 FILLER_35_1052 ();
 FILLCELL_X1 FILLER_35_1116 ();
 FILLCELL_X2 FILLER_35_1121 ();
 FILLCELL_X1 FILLER_35_1123 ();
 FILLCELL_X1 FILLER_35_1149 ();
 FILLCELL_X1 FILLER_35_1176 ();
 FILLCELL_X1 FILLER_35_1203 ();
 FILLCELL_X1 FILLER_35_1207 ();
 FILLCELL_X1 FILLER_35_1234 ();
 FILLCELL_X1 FILLER_35_1254 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X8 FILLER_36_97 ();
 FILLCELL_X2 FILLER_36_105 ();
 FILLCELL_X1 FILLER_36_107 ();
 FILLCELL_X2 FILLER_36_128 ();
 FILLCELL_X8 FILLER_36_164 ();
 FILLCELL_X4 FILLER_36_172 ();
 FILLCELL_X1 FILLER_36_176 ();
 FILLCELL_X4 FILLER_36_219 ();
 FILLCELL_X2 FILLER_36_223 ();
 FILLCELL_X1 FILLER_36_229 ();
 FILLCELL_X1 FILLER_36_234 ();
 FILLCELL_X8 FILLER_36_238 ();
 FILLCELL_X2 FILLER_36_246 ();
 FILLCELL_X4 FILLER_36_331 ();
 FILLCELL_X2 FILLER_36_335 ();
 FILLCELL_X1 FILLER_36_344 ();
 FILLCELL_X1 FILLER_36_359 ();
 FILLCELL_X8 FILLER_36_376 ();
 FILLCELL_X4 FILLER_36_384 ();
 FILLCELL_X2 FILLER_36_388 ();
 FILLCELL_X4 FILLER_36_397 ();
 FILLCELL_X2 FILLER_36_401 ();
 FILLCELL_X8 FILLER_36_406 ();
 FILLCELL_X4 FILLER_36_414 ();
 FILLCELL_X2 FILLER_36_418 ();
 FILLCELL_X1 FILLER_36_420 ();
 FILLCELL_X4 FILLER_36_441 ();
 FILLCELL_X1 FILLER_36_454 ();
 FILLCELL_X1 FILLER_36_462 ();
 FILLCELL_X1 FILLER_36_467 ();
 FILLCELL_X1 FILLER_36_475 ();
 FILLCELL_X1 FILLER_36_485 ();
 FILLCELL_X1 FILLER_36_493 ();
 FILLCELL_X4 FILLER_36_497 ();
 FILLCELL_X2 FILLER_36_531 ();
 FILLCELL_X1 FILLER_36_533 ();
 FILLCELL_X8 FILLER_36_541 ();
 FILLCELL_X1 FILLER_36_549 ();
 FILLCELL_X4 FILLER_36_570 ();
 FILLCELL_X1 FILLER_36_574 ();
 FILLCELL_X2 FILLER_36_604 ();
 FILLCELL_X1 FILLER_36_623 ();
 FILLCELL_X16 FILLER_36_632 ();
 FILLCELL_X8 FILLER_36_648 ();
 FILLCELL_X4 FILLER_36_730 ();
 FILLCELL_X16 FILLER_36_758 ();
 FILLCELL_X8 FILLER_36_774 ();
 FILLCELL_X4 FILLER_36_782 ();
 FILLCELL_X2 FILLER_36_786 ();
 FILLCELL_X2 FILLER_36_795 ();
 FILLCELL_X2 FILLER_36_812 ();
 FILLCELL_X4 FILLER_36_824 ();
 FILLCELL_X1 FILLER_36_828 ();
 FILLCELL_X8 FILLER_36_834 ();
 FILLCELL_X4 FILLER_36_842 ();
 FILLCELL_X2 FILLER_36_851 ();
 FILLCELL_X2 FILLER_36_860 ();
 FILLCELL_X4 FILLER_36_875 ();
 FILLCELL_X8 FILLER_36_888 ();
 FILLCELL_X1 FILLER_36_896 ();
 FILLCELL_X16 FILLER_36_908 ();
 FILLCELL_X8 FILLER_36_924 ();
 FILLCELL_X2 FILLER_36_932 ();
 FILLCELL_X4 FILLER_36_943 ();
 FILLCELL_X2 FILLER_36_964 ();
 FILLCELL_X2 FILLER_36_978 ();
 FILLCELL_X4 FILLER_36_1014 ();
 FILLCELL_X2 FILLER_36_1018 ();
 FILLCELL_X1 FILLER_36_1020 ();
 FILLCELL_X16 FILLER_36_1035 ();
 FILLCELL_X8 FILLER_36_1051 ();
 FILLCELL_X1 FILLER_36_1059 ();
 FILLCELL_X32 FILLER_36_1067 ();
 FILLCELL_X2 FILLER_36_1099 ();
 FILLCELL_X2 FILLER_36_1112 ();
 FILLCELL_X1 FILLER_36_1114 ();
 FILLCELL_X4 FILLER_36_1122 ();
 FILLCELL_X2 FILLER_36_1126 ();
 FILLCELL_X16 FILLER_36_1130 ();
 FILLCELL_X2 FILLER_36_1146 ();
 FILLCELL_X1 FILLER_36_1148 ();
 FILLCELL_X16 FILLER_36_1188 ();
 FILLCELL_X2 FILLER_36_1204 ();
 FILLCELL_X1 FILLER_36_1206 ();
 FILLCELL_X16 FILLER_36_1210 ();
 FILLCELL_X2 FILLER_36_1226 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X16 FILLER_37_65 ();
 FILLCELL_X4 FILLER_37_81 ();
 FILLCELL_X4 FILLER_37_152 ();
 FILLCELL_X2 FILLER_37_156 ();
 FILLCELL_X1 FILLER_37_158 ();
 FILLCELL_X1 FILLER_37_186 ();
 FILLCELL_X1 FILLER_37_201 ();
 FILLCELL_X4 FILLER_37_265 ();
 FILLCELL_X2 FILLER_37_269 ();
 FILLCELL_X1 FILLER_37_276 ();
 FILLCELL_X4 FILLER_37_280 ();
 FILLCELL_X1 FILLER_37_284 ();
 FILLCELL_X2 FILLER_37_289 ();
 FILLCELL_X2 FILLER_37_294 ();
 FILLCELL_X1 FILLER_37_296 ();
 FILLCELL_X8 FILLER_37_311 ();
 FILLCELL_X4 FILLER_37_319 ();
 FILLCELL_X1 FILLER_37_323 ();
 FILLCELL_X1 FILLER_37_331 ();
 FILLCELL_X1 FILLER_37_336 ();
 FILLCELL_X8 FILLER_37_340 ();
 FILLCELL_X1 FILLER_37_353 ();
 FILLCELL_X2 FILLER_37_357 ();
 FILLCELL_X1 FILLER_37_379 ();
 FILLCELL_X1 FILLER_37_404 ();
 FILLCELL_X1 FILLER_37_408 ();
 FILLCELL_X16 FILLER_37_429 ();
 FILLCELL_X4 FILLER_37_445 ();
 FILLCELL_X2 FILLER_37_449 ();
 FILLCELL_X1 FILLER_37_451 ();
 FILLCELL_X4 FILLER_37_470 ();
 FILLCELL_X1 FILLER_37_474 ();
 FILLCELL_X2 FILLER_37_490 ();
 FILLCELL_X8 FILLER_37_496 ();
 FILLCELL_X2 FILLER_37_504 ();
 FILLCELL_X8 FILLER_37_516 ();
 FILLCELL_X4 FILLER_37_524 ();
 FILLCELL_X2 FILLER_37_528 ();
 FILLCELL_X1 FILLER_37_544 ();
 FILLCELL_X8 FILLER_37_552 ();
 FILLCELL_X4 FILLER_37_591 ();
 FILLCELL_X1 FILLER_37_595 ();
 FILLCELL_X2 FILLER_37_605 ();
 FILLCELL_X4 FILLER_37_645 ();
 FILLCELL_X2 FILLER_37_658 ();
 FILLCELL_X1 FILLER_37_693 ();
 FILLCELL_X1 FILLER_37_698 ();
 FILLCELL_X1 FILLER_37_702 ();
 FILLCELL_X1 FILLER_37_710 ();
 FILLCELL_X1 FILLER_37_715 ();
 FILLCELL_X4 FILLER_37_721 ();
 FILLCELL_X1 FILLER_37_725 ();
 FILLCELL_X8 FILLER_37_737 ();
 FILLCELL_X1 FILLER_37_745 ();
 FILLCELL_X8 FILLER_37_760 ();
 FILLCELL_X4 FILLER_37_768 ();
 FILLCELL_X2 FILLER_37_772 ();
 FILLCELL_X4 FILLER_37_786 ();
 FILLCELL_X1 FILLER_37_812 ();
 FILLCELL_X4 FILLER_37_820 ();
 FILLCELL_X1 FILLER_37_824 ();
 FILLCELL_X1 FILLER_37_849 ();
 FILLCELL_X1 FILLER_37_854 ();
 FILLCELL_X2 FILLER_37_865 ();
 FILLCELL_X1 FILLER_37_871 ();
 FILLCELL_X4 FILLER_37_885 ();
 FILLCELL_X1 FILLER_37_889 ();
 FILLCELL_X1 FILLER_37_896 ();
 FILLCELL_X8 FILLER_37_900 ();
 FILLCELL_X1 FILLER_37_908 ();
 FILLCELL_X1 FILLER_37_916 ();
 FILLCELL_X8 FILLER_37_935 ();
 FILLCELL_X4 FILLER_37_943 ();
 FILLCELL_X2 FILLER_37_947 ();
 FILLCELL_X1 FILLER_37_949 ();
 FILLCELL_X2 FILLER_37_959 ();
 FILLCELL_X1 FILLER_37_961 ();
 FILLCELL_X2 FILLER_37_979 ();
 FILLCELL_X8 FILLER_37_986 ();
 FILLCELL_X4 FILLER_37_994 ();
 FILLCELL_X2 FILLER_37_998 ();
 FILLCELL_X1 FILLER_37_1000 ();
 FILLCELL_X4 FILLER_37_1008 ();
 FILLCELL_X1 FILLER_37_1012 ();
 FILLCELL_X16 FILLER_37_1033 ();
 FILLCELL_X8 FILLER_37_1049 ();
 FILLCELL_X1 FILLER_37_1057 ();
 FILLCELL_X2 FILLER_37_1072 ();
 FILLCELL_X1 FILLER_37_1074 ();
 FILLCELL_X4 FILLER_37_1082 ();
 FILLCELL_X2 FILLER_37_1086 ();
 FILLCELL_X1 FILLER_37_1088 ();
 FILLCELL_X4 FILLER_37_1094 ();
 FILLCELL_X1 FILLER_37_1114 ();
 FILLCELL_X1 FILLER_37_1124 ();
 FILLCELL_X1 FILLER_37_1143 ();
 FILLCELL_X2 FILLER_37_1168 ();
 FILLCELL_X1 FILLER_37_1170 ();
 FILLCELL_X2 FILLER_37_1198 ();
 FILLCELL_X2 FILLER_37_1207 ();
 FILLCELL_X1 FILLER_37_1209 ();
 FILLCELL_X1 FILLER_37_1224 ();
 FILLCELL_X2 FILLER_37_1228 ();
 FILLCELL_X1 FILLER_37_1230 ();
 FILLCELL_X2 FILLER_37_1238 ();
 FILLCELL_X2 FILLER_37_1247 ();
 FILLCELL_X2 FILLER_37_1253 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X16 FILLER_38_65 ();
 FILLCELL_X4 FILLER_38_81 ();
 FILLCELL_X2 FILLER_38_85 ();
 FILLCELL_X8 FILLER_38_94 ();
 FILLCELL_X2 FILLER_38_102 ();
 FILLCELL_X1 FILLER_38_104 ();
 FILLCELL_X8 FILLER_38_112 ();
 FILLCELL_X1 FILLER_38_135 ();
 FILLCELL_X4 FILLER_38_177 ();
 FILLCELL_X2 FILLER_38_181 ();
 FILLCELL_X4 FILLER_38_197 ();
 FILLCELL_X8 FILLER_38_215 ();
 FILLCELL_X4 FILLER_38_223 ();
 FILLCELL_X1 FILLER_38_227 ();
 FILLCELL_X16 FILLER_38_231 ();
 FILLCELL_X1 FILLER_38_247 ();
 FILLCELL_X2 FILLER_38_259 ();
 FILLCELL_X2 FILLER_38_268 ();
 FILLCELL_X1 FILLER_38_270 ();
 FILLCELL_X1 FILLER_38_311 ();
 FILLCELL_X2 FILLER_38_352 ();
 FILLCELL_X8 FILLER_38_381 ();
 FILLCELL_X2 FILLER_38_389 ();
 FILLCELL_X4 FILLER_38_398 ();
 FILLCELL_X16 FILLER_38_414 ();
 FILLCELL_X4 FILLER_38_430 ();
 FILLCELL_X4 FILLER_38_441 ();
 FILLCELL_X2 FILLER_38_445 ();
 FILLCELL_X1 FILLER_38_447 ();
 FILLCELL_X4 FILLER_38_474 ();
 FILLCELL_X1 FILLER_38_478 ();
 FILLCELL_X2 FILLER_38_495 ();
 FILLCELL_X1 FILLER_38_497 ();
 FILLCELL_X4 FILLER_38_503 ();
 FILLCELL_X1 FILLER_38_529 ();
 FILLCELL_X1 FILLER_38_533 ();
 FILLCELL_X1 FILLER_38_537 ();
 FILLCELL_X4 FILLER_38_542 ();
 FILLCELL_X2 FILLER_38_546 ();
 FILLCELL_X8 FILLER_38_555 ();
 FILLCELL_X2 FILLER_38_563 ();
 FILLCELL_X1 FILLER_38_565 ();
 FILLCELL_X8 FILLER_38_622 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X4 FILLER_38_639 ();
 FILLCELL_X1 FILLER_38_643 ();
 FILLCELL_X4 FILLER_38_674 ();
 FILLCELL_X2 FILLER_38_678 ();
 FILLCELL_X8 FILLER_38_703 ();
 FILLCELL_X4 FILLER_38_711 ();
 FILLCELL_X2 FILLER_38_715 ();
 FILLCELL_X4 FILLER_38_743 ();
 FILLCELL_X1 FILLER_38_747 ();
 FILLCELL_X4 FILLER_38_770 ();
 FILLCELL_X16 FILLER_38_794 ();
 FILLCELL_X4 FILLER_38_810 ();
 FILLCELL_X2 FILLER_38_814 ();
 FILLCELL_X1 FILLER_38_816 ();
 FILLCELL_X2 FILLER_38_824 ();
 FILLCELL_X8 FILLER_38_832 ();
 FILLCELL_X4 FILLER_38_840 ();
 FILLCELL_X4 FILLER_38_866 ();
 FILLCELL_X2 FILLER_38_870 ();
 FILLCELL_X1 FILLER_38_872 ();
 FILLCELL_X4 FILLER_38_908 ();
 FILLCELL_X2 FILLER_38_912 ();
 FILLCELL_X1 FILLER_38_914 ();
 FILLCELL_X8 FILLER_38_941 ();
 FILLCELL_X4 FILLER_38_949 ();
 FILLCELL_X1 FILLER_38_953 ();
 FILLCELL_X4 FILLER_38_963 ();
 FILLCELL_X2 FILLER_38_967 ();
 FILLCELL_X1 FILLER_38_969 ();
 FILLCELL_X1 FILLER_38_975 ();
 FILLCELL_X1 FILLER_38_981 ();
 FILLCELL_X1 FILLER_38_988 ();
 FILLCELL_X2 FILLER_38_1009 ();
 FILLCELL_X8 FILLER_38_1021 ();
 FILLCELL_X2 FILLER_38_1029 ();
 FILLCELL_X1 FILLER_38_1045 ();
 FILLCELL_X4 FILLER_38_1060 ();
 FILLCELL_X1 FILLER_38_1064 ();
 FILLCELL_X8 FILLER_38_1070 ();
 FILLCELL_X4 FILLER_38_1098 ();
 FILLCELL_X1 FILLER_38_1118 ();
 FILLCELL_X8 FILLER_38_1126 ();
 FILLCELL_X4 FILLER_38_1134 ();
 FILLCELL_X16 FILLER_38_1142 ();
 FILLCELL_X8 FILLER_38_1158 ();
 FILLCELL_X4 FILLER_38_1166 ();
 FILLCELL_X16 FILLER_38_1177 ();
 FILLCELL_X4 FILLER_38_1193 ();
 FILLCELL_X4 FILLER_38_1204 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X1 FILLER_39_65 ();
 FILLCELL_X16 FILLER_39_93 ();
 FILLCELL_X8 FILLER_39_109 ();
 FILLCELL_X4 FILLER_39_152 ();
 FILLCELL_X2 FILLER_39_156 ();
 FILLCELL_X1 FILLER_39_158 ();
 FILLCELL_X2 FILLER_39_164 ();
 FILLCELL_X2 FILLER_39_235 ();
 FILLCELL_X2 FILLER_39_241 ();
 FILLCELL_X1 FILLER_39_243 ();
 FILLCELL_X1 FILLER_39_267 ();
 FILLCELL_X2 FILLER_39_282 ();
 FILLCELL_X1 FILLER_39_284 ();
 FILLCELL_X2 FILLER_39_315 ();
 FILLCELL_X1 FILLER_39_317 ();
 FILLCELL_X1 FILLER_39_332 ();
 FILLCELL_X2 FILLER_39_337 ();
 FILLCELL_X4 FILLER_39_342 ();
 FILLCELL_X2 FILLER_39_346 ();
 FILLCELL_X1 FILLER_39_348 ();
 FILLCELL_X2 FILLER_39_418 ();
 FILLCELL_X16 FILLER_39_440 ();
 FILLCELL_X1 FILLER_39_456 ();
 FILLCELL_X2 FILLER_39_462 ();
 FILLCELL_X4 FILLER_39_485 ();
 FILLCELL_X4 FILLER_39_498 ();
 FILLCELL_X2 FILLER_39_502 ();
 FILLCELL_X2 FILLER_39_522 ();
 FILLCELL_X4 FILLER_39_548 ();
 FILLCELL_X2 FILLER_39_552 ();
 FILLCELL_X1 FILLER_39_554 ();
 FILLCELL_X8 FILLER_39_575 ();
 FILLCELL_X4 FILLER_39_583 ();
 FILLCELL_X1 FILLER_39_587 ();
 FILLCELL_X1 FILLER_39_595 ();
 FILLCELL_X4 FILLER_39_627 ();
 FILLCELL_X2 FILLER_39_631 ();
 FILLCELL_X1 FILLER_39_649 ();
 FILLCELL_X2 FILLER_39_662 ();
 FILLCELL_X1 FILLER_39_664 ();
 FILLCELL_X2 FILLER_39_672 ();
 FILLCELL_X1 FILLER_39_674 ();
 FILLCELL_X2 FILLER_39_685 ();
 FILLCELL_X2 FILLER_39_700 ();
 FILLCELL_X16 FILLER_39_708 ();
 FILLCELL_X4 FILLER_39_724 ();
 FILLCELL_X1 FILLER_39_728 ();
 FILLCELL_X2 FILLER_39_736 ();
 FILLCELL_X1 FILLER_39_738 ();
 FILLCELL_X2 FILLER_39_759 ();
 FILLCELL_X1 FILLER_39_761 ();
 FILLCELL_X8 FILLER_39_769 ();
 FILLCELL_X2 FILLER_39_777 ();
 FILLCELL_X1 FILLER_39_779 ();
 FILLCELL_X1 FILLER_39_782 ();
 FILLCELL_X2 FILLER_39_788 ();
 FILLCELL_X2 FILLER_39_802 ();
 FILLCELL_X1 FILLER_39_808 ();
 FILLCELL_X4 FILLER_39_816 ();
 FILLCELL_X1 FILLER_39_820 ();
 FILLCELL_X8 FILLER_39_831 ();
 FILLCELL_X4 FILLER_39_839 ();
 FILLCELL_X1 FILLER_39_843 ();
 FILLCELL_X4 FILLER_39_863 ();
 FILLCELL_X1 FILLER_39_875 ();
 FILLCELL_X2 FILLER_39_904 ();
 FILLCELL_X2 FILLER_39_927 ();
 FILLCELL_X1 FILLER_39_929 ();
 FILLCELL_X8 FILLER_39_952 ();
 FILLCELL_X4 FILLER_39_960 ();
 FILLCELL_X2 FILLER_39_964 ();
 FILLCELL_X1 FILLER_39_966 ();
 FILLCELL_X8 FILLER_39_969 ();
 FILLCELL_X8 FILLER_39_1016 ();
 FILLCELL_X4 FILLER_39_1024 ();
 FILLCELL_X2 FILLER_39_1028 ();
 FILLCELL_X4 FILLER_39_1083 ();
 FILLCELL_X1 FILLER_39_1114 ();
 FILLCELL_X1 FILLER_39_1120 ();
 FILLCELL_X1 FILLER_39_1141 ();
 FILLCELL_X8 FILLER_39_1147 ();
 FILLCELL_X2 FILLER_39_1155 ();
 FILLCELL_X4 FILLER_39_1204 ();
 FILLCELL_X1 FILLER_39_1254 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X16 FILLER_40_33 ();
 FILLCELL_X1 FILLER_40_49 ();
 FILLCELL_X1 FILLER_40_77 ();
 FILLCELL_X2 FILLER_40_139 ();
 FILLCELL_X1 FILLER_40_155 ();
 FILLCELL_X4 FILLER_40_183 ();
 FILLCELL_X2 FILLER_40_187 ();
 FILLCELL_X2 FILLER_40_196 ();
 FILLCELL_X1 FILLER_40_198 ();
 FILLCELL_X4 FILLER_40_322 ();
 FILLCELL_X1 FILLER_40_326 ();
 FILLCELL_X8 FILLER_40_347 ();
 FILLCELL_X2 FILLER_40_355 ();
 FILLCELL_X8 FILLER_40_382 ();
 FILLCELL_X4 FILLER_40_397 ();
 FILLCELL_X2 FILLER_40_401 ();
 FILLCELL_X1 FILLER_40_407 ();
 FILLCELL_X16 FILLER_40_411 ();
 FILLCELL_X8 FILLER_40_427 ();
 FILLCELL_X1 FILLER_40_442 ();
 FILLCELL_X4 FILLER_40_451 ();
 FILLCELL_X2 FILLER_40_458 ();
 FILLCELL_X8 FILLER_40_464 ();
 FILLCELL_X2 FILLER_40_472 ();
 FILLCELL_X1 FILLER_40_474 ();
 FILLCELL_X16 FILLER_40_480 ();
 FILLCELL_X2 FILLER_40_515 ();
 FILLCELL_X2 FILLER_40_526 ();
 FILLCELL_X2 FILLER_40_546 ();
 FILLCELL_X2 FILLER_40_555 ();
 FILLCELL_X1 FILLER_40_557 ();
 FILLCELL_X2 FILLER_40_565 ();
 FILLCELL_X1 FILLER_40_574 ();
 FILLCELL_X4 FILLER_40_582 ();
 FILLCELL_X2 FILLER_40_586 ();
 FILLCELL_X1 FILLER_40_588 ();
 FILLCELL_X2 FILLER_40_614 ();
 FILLCELL_X1 FILLER_40_616 ();
 FILLCELL_X4 FILLER_40_624 ();
 FILLCELL_X2 FILLER_40_628 ();
 FILLCELL_X1 FILLER_40_630 ();
 FILLCELL_X16 FILLER_40_662 ();
 FILLCELL_X8 FILLER_40_678 ();
 FILLCELL_X2 FILLER_40_686 ();
 FILLCELL_X1 FILLER_40_695 ();
 FILLCELL_X8 FILLER_40_702 ();
 FILLCELL_X4 FILLER_40_710 ();
 FILLCELL_X1 FILLER_40_714 ();
 FILLCELL_X1 FILLER_40_722 ();
 FILLCELL_X4 FILLER_40_730 ();
 FILLCELL_X2 FILLER_40_734 ();
 FILLCELL_X1 FILLER_40_736 ();
 FILLCELL_X1 FILLER_40_746 ();
 FILLCELL_X2 FILLER_40_751 ();
 FILLCELL_X1 FILLER_40_758 ();
 FILLCELL_X16 FILLER_40_773 ();
 FILLCELL_X2 FILLER_40_789 ();
 FILLCELL_X1 FILLER_40_791 ();
 FILLCELL_X4 FILLER_40_801 ();
 FILLCELL_X2 FILLER_40_844 ();
 FILLCELL_X1 FILLER_40_846 ();
 FILLCELL_X2 FILLER_40_863 ();
 FILLCELL_X8 FILLER_40_874 ();
 FILLCELL_X1 FILLER_40_882 ();
 FILLCELL_X2 FILLER_40_896 ();
 FILLCELL_X1 FILLER_40_898 ();
 FILLCELL_X2 FILLER_40_904 ();
 FILLCELL_X1 FILLER_40_906 ();
 FILLCELL_X2 FILLER_40_916 ();
 FILLCELL_X8 FILLER_40_940 ();
 FILLCELL_X1 FILLER_40_948 ();
 FILLCELL_X2 FILLER_40_963 ();
 FILLCELL_X1 FILLER_40_1014 ();
 FILLCELL_X2 FILLER_40_1035 ();
 FILLCELL_X2 FILLER_40_1044 ();
 FILLCELL_X2 FILLER_40_1053 ();
 FILLCELL_X4 FILLER_40_1062 ();
 FILLCELL_X4 FILLER_40_1072 ();
 FILLCELL_X4 FILLER_40_1081 ();
 FILLCELL_X8 FILLER_40_1103 ();
 FILLCELL_X4 FILLER_40_1111 ();
 FILLCELL_X8 FILLER_40_1121 ();
 FILLCELL_X4 FILLER_40_1129 ();
 FILLCELL_X2 FILLER_40_1133 ();
 FILLCELL_X1 FILLER_40_1152 ();
 FILLCELL_X8 FILLER_40_1206 ();
 FILLCELL_X1 FILLER_40_1214 ();
 FILLCELL_X1 FILLER_40_1242 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X16 FILLER_41_33 ();
 FILLCELL_X4 FILLER_41_49 ();
 FILLCELL_X1 FILLER_41_86 ();
 FILLCELL_X1 FILLER_41_94 ();
 FILLCELL_X4 FILLER_41_102 ();
 FILLCELL_X2 FILLER_41_106 ();
 FILLCELL_X1 FILLER_41_108 ();
 FILLCELL_X16 FILLER_41_120 ();
 FILLCELL_X8 FILLER_41_136 ();
 FILLCELL_X2 FILLER_41_144 ();
 FILLCELL_X4 FILLER_41_153 ();
 FILLCELL_X2 FILLER_41_157 ();
 FILLCELL_X1 FILLER_41_159 ();
 FILLCELL_X2 FILLER_41_180 ();
 FILLCELL_X1 FILLER_41_189 ();
 FILLCELL_X2 FILLER_41_204 ();
 FILLCELL_X1 FILLER_41_206 ();
 FILLCELL_X1 FILLER_41_224 ();
 FILLCELL_X2 FILLER_41_232 ();
 FILLCELL_X2 FILLER_41_254 ();
 FILLCELL_X1 FILLER_41_260 ();
 FILLCELL_X4 FILLER_41_271 ();
 FILLCELL_X2 FILLER_41_275 ();
 FILLCELL_X1 FILLER_41_277 ();
 FILLCELL_X16 FILLER_41_338 ();
 FILLCELL_X2 FILLER_41_354 ();
 FILLCELL_X4 FILLER_41_421 ();
 FILLCELL_X4 FILLER_41_445 ();
 FILLCELL_X4 FILLER_41_464 ();
 FILLCELL_X1 FILLER_41_468 ();
 FILLCELL_X8 FILLER_41_474 ();
 FILLCELL_X4 FILLER_41_482 ();
 FILLCELL_X2 FILLER_41_506 ();
 FILLCELL_X4 FILLER_41_514 ();
 FILLCELL_X2 FILLER_41_518 ();
 FILLCELL_X1 FILLER_41_520 ();
 FILLCELL_X2 FILLER_41_530 ();
 FILLCELL_X1 FILLER_41_532 ();
 FILLCELL_X8 FILLER_41_558 ();
 FILLCELL_X4 FILLER_41_566 ();
 FILLCELL_X2 FILLER_41_570 ();
 FILLCELL_X2 FILLER_41_576 ();
 FILLCELL_X1 FILLER_41_595 ();
 FILLCELL_X8 FILLER_41_631 ();
 FILLCELL_X2 FILLER_41_639 ();
 FILLCELL_X1 FILLER_41_641 ();
 FILLCELL_X1 FILLER_41_697 ();
 FILLCELL_X8 FILLER_41_719 ();
 FILLCELL_X4 FILLER_41_727 ();
 FILLCELL_X2 FILLER_41_763 ();
 FILLCELL_X1 FILLER_41_765 ();
 FILLCELL_X8 FILLER_41_831 ();
 FILLCELL_X1 FILLER_41_846 ();
 FILLCELL_X2 FILLER_41_854 ();
 FILLCELL_X1 FILLER_41_856 ();
 FILLCELL_X4 FILLER_41_866 ();
 FILLCELL_X1 FILLER_41_883 ();
 FILLCELL_X8 FILLER_41_893 ();
 FILLCELL_X2 FILLER_41_901 ();
 FILLCELL_X1 FILLER_41_903 ();
 FILLCELL_X4 FILLER_41_911 ();
 FILLCELL_X2 FILLER_41_915 ();
 FILLCELL_X1 FILLER_41_917 ();
 FILLCELL_X4 FILLER_41_927 ();
 FILLCELL_X4 FILLER_41_938 ();
 FILLCELL_X2 FILLER_41_942 ();
 FILLCELL_X8 FILLER_41_949 ();
 FILLCELL_X2 FILLER_41_957 ();
 FILLCELL_X1 FILLER_41_959 ();
 FILLCELL_X1 FILLER_41_972 ();
 FILLCELL_X4 FILLER_41_975 ();
 FILLCELL_X1 FILLER_41_979 ();
 FILLCELL_X8 FILLER_41_987 ();
 FILLCELL_X1 FILLER_41_1007 ();
 FILLCELL_X16 FILLER_41_1012 ();
 FILLCELL_X8 FILLER_41_1028 ();
 FILLCELL_X4 FILLER_41_1036 ();
 FILLCELL_X4 FILLER_41_1054 ();
 FILLCELL_X8 FILLER_41_1078 ();
 FILLCELL_X1 FILLER_41_1086 ();
 FILLCELL_X1 FILLER_41_1110 ();
 FILLCELL_X2 FILLER_41_1126 ();
 FILLCELL_X4 FILLER_41_1144 ();
 FILLCELL_X4 FILLER_41_1153 ();
 FILLCELL_X1 FILLER_41_1157 ();
 FILLCELL_X1 FILLER_41_1192 ();
 FILLCELL_X8 FILLER_41_1220 ();
 FILLCELL_X2 FILLER_41_1228 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X8 FILLER_42_33 ();
 FILLCELL_X4 FILLER_42_41 ();
 FILLCELL_X1 FILLER_42_45 ();
 FILLCELL_X4 FILLER_42_88 ();
 FILLCELL_X1 FILLER_42_157 ();
 FILLCELL_X1 FILLER_42_165 ();
 FILLCELL_X4 FILLER_42_173 ();
 FILLCELL_X1 FILLER_42_177 ();
 FILLCELL_X1 FILLER_42_205 ();
 FILLCELL_X2 FILLER_42_227 ();
 FILLCELL_X8 FILLER_42_269 ();
 FILLCELL_X1 FILLER_42_277 ();
 FILLCELL_X1 FILLER_42_303 ();
 FILLCELL_X1 FILLER_42_311 ();
 FILLCELL_X4 FILLER_42_339 ();
 FILLCELL_X4 FILLER_42_347 ();
 FILLCELL_X8 FILLER_42_354 ();
 FILLCELL_X2 FILLER_42_382 ();
 FILLCELL_X4 FILLER_42_388 ();
 FILLCELL_X2 FILLER_42_392 ();
 FILLCELL_X1 FILLER_42_394 ();
 FILLCELL_X8 FILLER_42_415 ();
 FILLCELL_X4 FILLER_42_428 ();
 FILLCELL_X1 FILLER_42_439 ();
 FILLCELL_X2 FILLER_42_447 ();
 FILLCELL_X1 FILLER_42_456 ();
 FILLCELL_X2 FILLER_42_461 ();
 FILLCELL_X2 FILLER_42_467 ();
 FILLCELL_X1 FILLER_42_469 ();
 FILLCELL_X4 FILLER_42_484 ();
 FILLCELL_X2 FILLER_42_488 ();
 FILLCELL_X2 FILLER_42_524 ();
 FILLCELL_X1 FILLER_42_526 ();
 FILLCELL_X1 FILLER_42_532 ();
 FILLCELL_X1 FILLER_42_537 ();
 FILLCELL_X8 FILLER_42_547 ();
 FILLCELL_X1 FILLER_42_555 ();
 FILLCELL_X16 FILLER_42_560 ();
 FILLCELL_X8 FILLER_42_576 ();
 FILLCELL_X4 FILLER_42_584 ();
 FILLCELL_X2 FILLER_42_592 ();
 FILLCELL_X1 FILLER_42_594 ();
 FILLCELL_X16 FILLER_42_598 ();
 FILLCELL_X8 FILLER_42_614 ();
 FILLCELL_X4 FILLER_42_626 ();
 FILLCELL_X1 FILLER_42_630 ();
 FILLCELL_X4 FILLER_42_677 ();
 FILLCELL_X2 FILLER_42_698 ();
 FILLCELL_X1 FILLER_42_700 ();
 FILLCELL_X2 FILLER_42_730 ();
 FILLCELL_X1 FILLER_42_732 ();
 FILLCELL_X1 FILLER_42_762 ();
 FILLCELL_X8 FILLER_42_775 ();
 FILLCELL_X2 FILLER_42_783 ();
 FILLCELL_X1 FILLER_42_785 ();
 FILLCELL_X2 FILLER_42_793 ();
 FILLCELL_X4 FILLER_42_809 ();
 FILLCELL_X2 FILLER_42_813 ();
 FILLCELL_X1 FILLER_42_826 ();
 FILLCELL_X4 FILLER_42_832 ();
 FILLCELL_X2 FILLER_42_836 ();
 FILLCELL_X1 FILLER_42_838 ();
 FILLCELL_X4 FILLER_42_855 ();
 FILLCELL_X2 FILLER_42_859 ();
 FILLCELL_X1 FILLER_42_861 ();
 FILLCELL_X2 FILLER_42_873 ();
 FILLCELL_X2 FILLER_42_884 ();
 FILLCELL_X1 FILLER_42_886 ();
 FILLCELL_X1 FILLER_42_905 ();
 FILLCELL_X2 FILLER_42_915 ();
 FILLCELL_X1 FILLER_42_917 ();
 FILLCELL_X16 FILLER_42_927 ();
 FILLCELL_X1 FILLER_42_965 ();
 FILLCELL_X1 FILLER_42_970 ();
 FILLCELL_X8 FILLER_42_994 ();
 FILLCELL_X4 FILLER_42_1002 ();
 FILLCELL_X2 FILLER_42_1006 ();
 FILLCELL_X1 FILLER_42_1008 ();
 FILLCELL_X1 FILLER_42_1029 ();
 FILLCELL_X2 FILLER_42_1034 ();
 FILLCELL_X4 FILLER_42_1056 ();
 FILLCELL_X1 FILLER_42_1065 ();
 FILLCELL_X2 FILLER_42_1068 ();
 FILLCELL_X2 FILLER_42_1083 ();
 FILLCELL_X1 FILLER_42_1085 ();
 FILLCELL_X4 FILLER_42_1090 ();
 FILLCELL_X1 FILLER_42_1094 ();
 FILLCELL_X4 FILLER_42_1098 ();
 FILLCELL_X1 FILLER_42_1102 ();
 FILLCELL_X2 FILLER_42_1110 ();
 FILLCELL_X2 FILLER_42_1117 ();
 FILLCELL_X8 FILLER_42_1126 ();
 FILLCELL_X4 FILLER_42_1134 ();
 FILLCELL_X2 FILLER_42_1156 ();
 FILLCELL_X1 FILLER_42_1158 ();
 FILLCELL_X1 FILLER_42_1162 ();
 FILLCELL_X1 FILLER_42_1174 ();
 FILLCELL_X1 FILLER_42_1200 ();
 FILLCELL_X2 FILLER_42_1249 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X16 FILLER_43_33 ();
 FILLCELL_X2 FILLER_43_56 ();
 FILLCELL_X1 FILLER_43_58 ();
 FILLCELL_X1 FILLER_43_93 ();
 FILLCELL_X4 FILLER_43_101 ();
 FILLCELL_X4 FILLER_43_112 ();
 FILLCELL_X1 FILLER_43_116 ();
 FILLCELL_X1 FILLER_43_138 ();
 FILLCELL_X2 FILLER_43_153 ();
 FILLCELL_X1 FILLER_43_211 ();
 FILLCELL_X2 FILLER_43_239 ();
 FILLCELL_X2 FILLER_43_252 ();
 FILLCELL_X4 FILLER_43_268 ();
 FILLCELL_X8 FILLER_43_286 ();
 FILLCELL_X4 FILLER_43_294 ();
 FILLCELL_X2 FILLER_43_298 ();
 FILLCELL_X2 FILLER_43_350 ();
 FILLCELL_X1 FILLER_43_352 ();
 FILLCELL_X8 FILLER_43_356 ();
 FILLCELL_X2 FILLER_43_364 ();
 FILLCELL_X2 FILLER_43_400 ();
 FILLCELL_X4 FILLER_43_408 ();
 FILLCELL_X2 FILLER_43_412 ();
 FILLCELL_X1 FILLER_43_414 ();
 FILLCELL_X4 FILLER_43_437 ();
 FILLCELL_X2 FILLER_43_450 ();
 FILLCELL_X2 FILLER_43_466 ();
 FILLCELL_X4 FILLER_43_473 ();
 FILLCELL_X4 FILLER_43_497 ();
 FILLCELL_X1 FILLER_43_501 ();
 FILLCELL_X8 FILLER_43_519 ();
 FILLCELL_X2 FILLER_43_527 ();
 FILLCELL_X4 FILLER_43_544 ();
 FILLCELL_X1 FILLER_43_548 ();
 FILLCELL_X2 FILLER_43_558 ();
 FILLCELL_X1 FILLER_43_560 ();
 FILLCELL_X4 FILLER_43_581 ();
 FILLCELL_X2 FILLER_43_602 ();
 FILLCELL_X1 FILLER_43_604 ();
 FILLCELL_X4 FILLER_43_622 ();
 FILLCELL_X1 FILLER_43_626 ();
 FILLCELL_X2 FILLER_43_636 ();
 FILLCELL_X2 FILLER_43_656 ();
 FILLCELL_X1 FILLER_43_658 ();
 FILLCELL_X2 FILLER_43_689 ();
 FILLCELL_X2 FILLER_43_694 ();
 FILLCELL_X16 FILLER_43_701 ();
 FILLCELL_X2 FILLER_43_717 ();
 FILLCELL_X1 FILLER_43_719 ();
 FILLCELL_X2 FILLER_43_739 ();
 FILLCELL_X1 FILLER_43_741 ();
 FILLCELL_X1 FILLER_43_747 ();
 FILLCELL_X1 FILLER_43_756 ();
 FILLCELL_X8 FILLER_43_787 ();
 FILLCELL_X1 FILLER_43_795 ();
 FILLCELL_X8 FILLER_43_802 ();
 FILLCELL_X4 FILLER_43_810 ();
 FILLCELL_X8 FILLER_43_831 ();
 FILLCELL_X4 FILLER_43_839 ();
 FILLCELL_X2 FILLER_43_852 ();
 FILLCELL_X1 FILLER_43_854 ();
 FILLCELL_X2 FILLER_43_859 ();
 FILLCELL_X1 FILLER_43_861 ();
 FILLCELL_X4 FILLER_43_870 ();
 FILLCELL_X1 FILLER_43_881 ();
 FILLCELL_X4 FILLER_43_891 ();
 FILLCELL_X2 FILLER_43_895 ();
 FILLCELL_X8 FILLER_43_904 ();
 FILLCELL_X1 FILLER_43_912 ();
 FILLCELL_X16 FILLER_43_930 ();
 FILLCELL_X4 FILLER_43_946 ();
 FILLCELL_X2 FILLER_43_950 ();
 FILLCELL_X8 FILLER_43_954 ();
 FILLCELL_X4 FILLER_43_962 ();
 FILLCELL_X2 FILLER_43_966 ();
 FILLCELL_X1 FILLER_43_979 ();
 FILLCELL_X2 FILLER_43_982 ();
 FILLCELL_X1 FILLER_43_984 ();
 FILLCELL_X2 FILLER_43_1012 ();
 FILLCELL_X1 FILLER_43_1014 ();
 FILLCELL_X4 FILLER_43_1022 ();
 FILLCELL_X2 FILLER_43_1026 ();
 FILLCELL_X2 FILLER_43_1042 ();
 FILLCELL_X1 FILLER_43_1044 ();
 FILLCELL_X2 FILLER_43_1052 ();
 FILLCELL_X1 FILLER_43_1054 ();
 FILLCELL_X8 FILLER_43_1065 ();
 FILLCELL_X4 FILLER_43_1073 ();
 FILLCELL_X2 FILLER_43_1077 ();
 FILLCELL_X2 FILLER_43_1102 ();
 FILLCELL_X8 FILLER_43_1124 ();
 FILLCELL_X2 FILLER_43_1132 ();
 FILLCELL_X2 FILLER_43_1142 ();
 FILLCELL_X1 FILLER_43_1144 ();
 FILLCELL_X4 FILLER_43_1149 ();
 FILLCELL_X2 FILLER_43_1153 ();
 FILLCELL_X1 FILLER_43_1155 ();
 FILLCELL_X8 FILLER_43_1167 ();
 FILLCELL_X2 FILLER_43_1175 ();
 FILLCELL_X8 FILLER_43_1186 ();
 FILLCELL_X4 FILLER_43_1194 ();
 FILLCELL_X2 FILLER_43_1198 ();
 FILLCELL_X1 FILLER_43_1200 ();
 FILLCELL_X1 FILLER_43_1212 ();
 FILLCELL_X8 FILLER_43_1219 ();
 FILLCELL_X1 FILLER_43_1230 ();
 FILLCELL_X1 FILLER_43_1239 ();
 FILLCELL_X2 FILLER_43_1244 ();
 FILLCELL_X1 FILLER_43_1246 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X2 FILLER_44_33 ();
 FILLCELL_X1 FILLER_44_35 ();
 FILLCELL_X1 FILLER_44_56 ();
 FILLCELL_X2 FILLER_44_64 ();
 FILLCELL_X1 FILLER_44_85 ();
 FILLCELL_X16 FILLER_44_93 ();
 FILLCELL_X2 FILLER_44_109 ();
 FILLCELL_X4 FILLER_44_131 ();
 FILLCELL_X2 FILLER_44_135 ();
 FILLCELL_X2 FILLER_44_225 ();
 FILLCELL_X16 FILLER_44_277 ();
 FILLCELL_X1 FILLER_44_293 ();
 FILLCELL_X4 FILLER_44_314 ();
 FILLCELL_X1 FILLER_44_318 ();
 FILLCELL_X1 FILLER_44_333 ();
 FILLCELL_X1 FILLER_44_388 ();
 FILLCELL_X1 FILLER_44_401 ();
 FILLCELL_X2 FILLER_44_422 ();
 FILLCELL_X2 FILLER_44_458 ();
 FILLCELL_X1 FILLER_44_460 ();
 FILLCELL_X2 FILLER_44_468 ();
 FILLCELL_X2 FILLER_44_482 ();
 FILLCELL_X4 FILLER_44_491 ();
 FILLCELL_X4 FILLER_44_499 ();
 FILLCELL_X2 FILLER_44_512 ();
 FILLCELL_X2 FILLER_44_516 ();
 FILLCELL_X2 FILLER_44_525 ();
 FILLCELL_X2 FILLER_44_555 ();
 FILLCELL_X1 FILLER_44_557 ();
 FILLCELL_X8 FILLER_44_582 ();
 FILLCELL_X8 FILLER_44_593 ();
 FILLCELL_X1 FILLER_44_601 ();
 FILLCELL_X4 FILLER_44_616 ();
 FILLCELL_X1 FILLER_44_620 ();
 FILLCELL_X1 FILLER_44_630 ();
 FILLCELL_X4 FILLER_44_639 ();
 FILLCELL_X1 FILLER_44_657 ();
 FILLCELL_X8 FILLER_44_679 ();
 FILLCELL_X4 FILLER_44_687 ();
 FILLCELL_X2 FILLER_44_691 ();
 FILLCELL_X1 FILLER_44_693 ();
 FILLCELL_X2 FILLER_44_721 ();
 FILLCELL_X1 FILLER_44_723 ();
 FILLCELL_X4 FILLER_44_741 ();
 FILLCELL_X1 FILLER_44_756 ();
 FILLCELL_X2 FILLER_44_777 ();
 FILLCELL_X1 FILLER_44_779 ();
 FILLCELL_X4 FILLER_44_805 ();
 FILLCELL_X4 FILLER_44_824 ();
 FILLCELL_X2 FILLER_44_828 ();
 FILLCELL_X2 FILLER_44_833 ();
 FILLCELL_X2 FILLER_44_844 ();
 FILLCELL_X1 FILLER_44_846 ();
 FILLCELL_X1 FILLER_44_852 ();
 FILLCELL_X2 FILLER_44_857 ();
 FILLCELL_X2 FILLER_44_877 ();
 FILLCELL_X8 FILLER_44_906 ();
 FILLCELL_X4 FILLER_44_914 ();
 FILLCELL_X2 FILLER_44_918 ();
 FILLCELL_X16 FILLER_44_929 ();
 FILLCELL_X4 FILLER_44_945 ();
 FILLCELL_X1 FILLER_44_951 ();
 FILLCELL_X1 FILLER_44_956 ();
 FILLCELL_X1 FILLER_44_961 ();
 FILLCELL_X1 FILLER_44_965 ();
 FILLCELL_X2 FILLER_44_975 ();
 FILLCELL_X16 FILLER_44_991 ();
 FILLCELL_X4 FILLER_44_1007 ();
 FILLCELL_X4 FILLER_44_1024 ();
 FILLCELL_X1 FILLER_44_1028 ();
 FILLCELL_X8 FILLER_44_1032 ();
 FILLCELL_X2 FILLER_44_1040 ();
 FILLCELL_X2 FILLER_44_1054 ();
 FILLCELL_X1 FILLER_44_1056 ();
 FILLCELL_X4 FILLER_44_1082 ();
 FILLCELL_X1 FILLER_44_1108 ();
 FILLCELL_X1 FILLER_44_1114 ();
 FILLCELL_X4 FILLER_44_1154 ();
 FILLCELL_X4 FILLER_44_1165 ();
 FILLCELL_X1 FILLER_44_1169 ();
 FILLCELL_X1 FILLER_44_1177 ();
 FILLCELL_X4 FILLER_44_1200 ();
 FILLCELL_X1 FILLER_44_1204 ();
 FILLCELL_X2 FILLER_44_1217 ();
 FILLCELL_X4 FILLER_44_1230 ();
 FILLCELL_X1 FILLER_44_1234 ();
 FILLCELL_X8 FILLER_44_1244 ();
 FILLCELL_X2 FILLER_44_1252 ();
 FILLCELL_X1 FILLER_44_1254 ();
 FILLCELL_X16 FILLER_45_1 ();
 FILLCELL_X4 FILLER_45_44 ();
 FILLCELL_X2 FILLER_45_48 ();
 FILLCELL_X2 FILLER_45_84 ();
 FILLCELL_X1 FILLER_45_86 ();
 FILLCELL_X2 FILLER_45_108 ();
 FILLCELL_X1 FILLER_45_110 ();
 FILLCELL_X16 FILLER_45_118 ();
 FILLCELL_X1 FILLER_45_255 ();
 FILLCELL_X1 FILLER_45_263 ();
 FILLCELL_X4 FILLER_45_342 ();
 FILLCELL_X4 FILLER_45_350 ();
 FILLCELL_X2 FILLER_45_354 ();
 FILLCELL_X2 FILLER_45_359 ();
 FILLCELL_X1 FILLER_45_361 ();
 FILLCELL_X4 FILLER_45_375 ();
 FILLCELL_X1 FILLER_45_379 ();
 FILLCELL_X16 FILLER_45_408 ();
 FILLCELL_X8 FILLER_45_424 ();
 FILLCELL_X4 FILLER_45_432 ();
 FILLCELL_X1 FILLER_45_436 ();
 FILLCELL_X1 FILLER_45_449 ();
 FILLCELL_X4 FILLER_45_457 ();
 FILLCELL_X1 FILLER_45_461 ();
 FILLCELL_X4 FILLER_45_487 ();
 FILLCELL_X8 FILLER_45_520 ();
 FILLCELL_X4 FILLER_45_528 ();
 FILLCELL_X2 FILLER_45_535 ();
 FILLCELL_X1 FILLER_45_537 ();
 FILLCELL_X4 FILLER_45_545 ();
 FILLCELL_X2 FILLER_45_549 ();
 FILLCELL_X4 FILLER_45_564 ();
 FILLCELL_X1 FILLER_45_568 ();
 FILLCELL_X16 FILLER_45_596 ();
 FILLCELL_X1 FILLER_45_612 ();
 FILLCELL_X4 FILLER_45_617 ();
 FILLCELL_X2 FILLER_45_621 ();
 FILLCELL_X1 FILLER_45_623 ();
 FILLCELL_X16 FILLER_45_682 ();
 FILLCELL_X2 FILLER_45_698 ();
 FILLCELL_X1 FILLER_45_700 ();
 FILLCELL_X4 FILLER_45_726 ();
 FILLCELL_X1 FILLER_45_730 ();
 FILLCELL_X1 FILLER_45_734 ();
 FILLCELL_X2 FILLER_45_739 ();
 FILLCELL_X1 FILLER_45_745 ();
 FILLCELL_X1 FILLER_45_750 ();
 FILLCELL_X16 FILLER_45_768 ();
 FILLCELL_X2 FILLER_45_784 ();
 FILLCELL_X2 FILLER_45_795 ();
 FILLCELL_X1 FILLER_45_797 ();
 FILLCELL_X1 FILLER_45_824 ();
 FILLCELL_X1 FILLER_45_834 ();
 FILLCELL_X2 FILLER_45_839 ();
 FILLCELL_X2 FILLER_45_844 ();
 FILLCELL_X2 FILLER_45_850 ();
 FILLCELL_X1 FILLER_45_856 ();
 FILLCELL_X4 FILLER_45_877 ();
 FILLCELL_X2 FILLER_45_881 ();
 FILLCELL_X16 FILLER_45_901 ();
 FILLCELL_X8 FILLER_45_917 ();
 FILLCELL_X4 FILLER_45_945 ();
 FILLCELL_X1 FILLER_45_957 ();
 FILLCELL_X8 FILLER_45_981 ();
 FILLCELL_X1 FILLER_45_989 ();
 FILLCELL_X2 FILLER_45_1002 ();
 FILLCELL_X2 FILLER_45_1100 ();
 FILLCELL_X1 FILLER_45_1102 ();
 FILLCELL_X16 FILLER_45_1105 ();
 FILLCELL_X2 FILLER_45_1121 ();
 FILLCELL_X2 FILLER_45_1133 ();
 FILLCELL_X1 FILLER_45_1135 ();
 FILLCELL_X2 FILLER_45_1143 ();
 FILLCELL_X4 FILLER_45_1165 ();
 FILLCELL_X4 FILLER_45_1189 ();
 FILLCELL_X2 FILLER_45_1213 ();
 FILLCELL_X1 FILLER_45_1215 ();
 FILLCELL_X4 FILLER_45_1220 ();
 FILLCELL_X2 FILLER_45_1224 ();
 FILLCELL_X1 FILLER_45_1226 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X8 FILLER_46_33 ();
 FILLCELL_X4 FILLER_46_41 ();
 FILLCELL_X2 FILLER_46_45 ();
 FILLCELL_X1 FILLER_46_47 ();
 FILLCELL_X2 FILLER_46_55 ();
 FILLCELL_X1 FILLER_46_57 ();
 FILLCELL_X1 FILLER_46_86 ();
 FILLCELL_X4 FILLER_46_114 ();
 FILLCELL_X2 FILLER_46_118 ();
 FILLCELL_X1 FILLER_46_120 ();
 FILLCELL_X1 FILLER_46_154 ();
 FILLCELL_X2 FILLER_46_250 ();
 FILLCELL_X4 FILLER_46_259 ();
 FILLCELL_X2 FILLER_46_263 ();
 FILLCELL_X8 FILLER_46_274 ();
 FILLCELL_X4 FILLER_46_282 ();
 FILLCELL_X2 FILLER_46_286 ();
 FILLCELL_X1 FILLER_46_288 ();
 FILLCELL_X8 FILLER_46_292 ();
 FILLCELL_X4 FILLER_46_300 ();
 FILLCELL_X2 FILLER_46_304 ();
 FILLCELL_X1 FILLER_46_306 ();
 FILLCELL_X4 FILLER_46_316 ();
 FILLCELL_X8 FILLER_46_327 ();
 FILLCELL_X2 FILLER_46_362 ();
 FILLCELL_X4 FILLER_46_377 ();
 FILLCELL_X2 FILLER_46_381 ();
 FILLCELL_X1 FILLER_46_390 ();
 FILLCELL_X2 FILLER_46_398 ();
 FILLCELL_X2 FILLER_46_407 ();
 FILLCELL_X4 FILLER_46_416 ();
 FILLCELL_X2 FILLER_46_440 ();
 FILLCELL_X4 FILLER_46_449 ();
 FILLCELL_X2 FILLER_46_453 ();
 FILLCELL_X1 FILLER_46_455 ();
 FILLCELL_X2 FILLER_46_459 ();
 FILLCELL_X1 FILLER_46_461 ();
 FILLCELL_X1 FILLER_46_469 ();
 FILLCELL_X2 FILLER_46_472 ();
 FILLCELL_X8 FILLER_46_481 ();
 FILLCELL_X1 FILLER_46_489 ();
 FILLCELL_X4 FILLER_46_504 ();
 FILLCELL_X2 FILLER_46_508 ();
 FILLCELL_X1 FILLER_46_526 ();
 FILLCELL_X2 FILLER_46_534 ();
 FILLCELL_X2 FILLER_46_539 ();
 FILLCELL_X2 FILLER_46_548 ();
 FILLCELL_X1 FILLER_46_550 ();
 FILLCELL_X8 FILLER_46_554 ();
 FILLCELL_X8 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_617 ();
 FILLCELL_X1 FILLER_46_621 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X4 FILLER_46_632 ();
 FILLCELL_X1 FILLER_46_649 ();
 FILLCELL_X4 FILLER_46_659 ();
 FILLCELL_X2 FILLER_46_663 ();
 FILLCELL_X1 FILLER_46_665 ();
 FILLCELL_X2 FILLER_46_702 ();
 FILLCELL_X1 FILLER_46_704 ();
 FILLCELL_X4 FILLER_46_714 ();
 FILLCELL_X2 FILLER_46_718 ();
 FILLCELL_X1 FILLER_46_720 ();
 FILLCELL_X2 FILLER_46_739 ();
 FILLCELL_X8 FILLER_46_746 ();
 FILLCELL_X4 FILLER_46_754 ();
 FILLCELL_X1 FILLER_46_758 ();
 FILLCELL_X16 FILLER_46_773 ();
 FILLCELL_X8 FILLER_46_789 ();
 FILLCELL_X4 FILLER_46_797 ();
 FILLCELL_X2 FILLER_46_801 ();
 FILLCELL_X1 FILLER_46_866 ();
 FILLCELL_X8 FILLER_46_873 ();
 FILLCELL_X4 FILLER_46_881 ();
 FILLCELL_X2 FILLER_46_904 ();
 FILLCELL_X1 FILLER_46_906 ();
 FILLCELL_X1 FILLER_46_932 ();
 FILLCELL_X2 FILLER_46_955 ();
 FILLCELL_X2 FILLER_46_961 ();
 FILLCELL_X4 FILLER_46_968 ();
 FILLCELL_X1 FILLER_46_972 ();
 FILLCELL_X2 FILLER_46_995 ();
 FILLCELL_X2 FILLER_46_1043 ();
 FILLCELL_X1 FILLER_46_1049 ();
 FILLCELL_X32 FILLER_46_1054 ();
 FILLCELL_X4 FILLER_46_1086 ();
 FILLCELL_X2 FILLER_46_1090 ();
 FILLCELL_X1 FILLER_46_1092 ();
 FILLCELL_X8 FILLER_46_1100 ();
 FILLCELL_X4 FILLER_46_1108 ();
 FILLCELL_X2 FILLER_46_1112 ();
 FILLCELL_X2 FILLER_46_1121 ();
 FILLCELL_X1 FILLER_46_1123 ();
 FILLCELL_X8 FILLER_46_1151 ();
 FILLCELL_X4 FILLER_46_1159 ();
 FILLCELL_X16 FILLER_46_1170 ();
 FILLCELL_X4 FILLER_46_1186 ();
 FILLCELL_X2 FILLER_46_1190 ();
 FILLCELL_X2 FILLER_46_1199 ();
 FILLCELL_X1 FILLER_46_1201 ();
 FILLCELL_X1 FILLER_46_1224 ();
 FILLCELL_X1 FILLER_46_1227 ();
 FILLCELL_X1 FILLER_46_1232 ();
 FILLCELL_X4 FILLER_46_1240 ();
 FILLCELL_X1 FILLER_46_1244 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X4 FILLER_47_17 ();
 FILLCELL_X1 FILLER_47_21 ();
 FILLCELL_X4 FILLER_47_29 ();
 FILLCELL_X2 FILLER_47_53 ();
 FILLCELL_X1 FILLER_47_55 ();
 FILLCELL_X4 FILLER_47_76 ();
 FILLCELL_X2 FILLER_47_80 ();
 FILLCELL_X2 FILLER_47_102 ();
 FILLCELL_X1 FILLER_47_104 ();
 FILLCELL_X4 FILLER_47_112 ();
 FILLCELL_X2 FILLER_47_116 ();
 FILLCELL_X4 FILLER_47_138 ();
 FILLCELL_X2 FILLER_47_142 ();
 FILLCELL_X2 FILLER_47_257 ();
 FILLCELL_X8 FILLER_47_269 ();
 FILLCELL_X2 FILLER_47_281 ();
 FILLCELL_X8 FILLER_47_303 ();
 FILLCELL_X2 FILLER_47_311 ();
 FILLCELL_X1 FILLER_47_313 ();
 FILLCELL_X4 FILLER_47_317 ();
 FILLCELL_X2 FILLER_47_335 ();
 FILLCELL_X2 FILLER_47_358 ();
 FILLCELL_X1 FILLER_47_360 ();
 FILLCELL_X16 FILLER_47_381 ();
 FILLCELL_X4 FILLER_47_397 ();
 FILLCELL_X8 FILLER_47_408 ();
 FILLCELL_X4 FILLER_47_420 ();
 FILLCELL_X1 FILLER_47_424 ();
 FILLCELL_X4 FILLER_47_428 ();
 FILLCELL_X2 FILLER_47_432 ();
 FILLCELL_X1 FILLER_47_434 ();
 FILLCELL_X4 FILLER_47_442 ();
 FILLCELL_X2 FILLER_47_470 ();
 FILLCELL_X8 FILLER_47_476 ();
 FILLCELL_X4 FILLER_47_484 ();
 FILLCELL_X1 FILLER_47_491 ();
 FILLCELL_X4 FILLER_47_503 ();
 FILLCELL_X2 FILLER_47_507 ();
 FILLCELL_X4 FILLER_47_522 ();
 FILLCELL_X8 FILLER_47_533 ();
 FILLCELL_X2 FILLER_47_541 ();
 FILLCELL_X1 FILLER_47_543 ();
 FILLCELL_X1 FILLER_47_572 ();
 FILLCELL_X4 FILLER_47_583 ();
 FILLCELL_X1 FILLER_47_587 ();
 FILLCELL_X1 FILLER_47_595 ();
 FILLCELL_X4 FILLER_47_629 ();
 FILLCELL_X2 FILLER_47_633 ();
 FILLCELL_X1 FILLER_47_635 ();
 FILLCELL_X1 FILLER_47_657 ();
 FILLCELL_X8 FILLER_47_670 ();
 FILLCELL_X4 FILLER_47_678 ();
 FILLCELL_X8 FILLER_47_693 ();
 FILLCELL_X2 FILLER_47_701 ();
 FILLCELL_X4 FILLER_47_723 ();
 FILLCELL_X2 FILLER_47_727 ();
 FILLCELL_X1 FILLER_47_729 ();
 FILLCELL_X1 FILLER_47_734 ();
 FILLCELL_X2 FILLER_47_747 ();
 FILLCELL_X1 FILLER_47_749 ();
 FILLCELL_X1 FILLER_47_761 ();
 FILLCELL_X16 FILLER_47_774 ();
 FILLCELL_X1 FILLER_47_790 ();
 FILLCELL_X8 FILLER_47_816 ();
 FILLCELL_X1 FILLER_47_824 ();
 FILLCELL_X8 FILLER_47_832 ();
 FILLCELL_X1 FILLER_47_843 ();
 FILLCELL_X1 FILLER_47_848 ();
 FILLCELL_X1 FILLER_47_856 ();
 FILLCELL_X2 FILLER_47_862 ();
 FILLCELL_X1 FILLER_47_864 ();
 FILLCELL_X4 FILLER_47_870 ();
 FILLCELL_X2 FILLER_47_874 ();
 FILLCELL_X1 FILLER_47_876 ();
 FILLCELL_X2 FILLER_47_895 ();
 FILLCELL_X1 FILLER_47_907 ();
 FILLCELL_X2 FILLER_47_912 ();
 FILLCELL_X1 FILLER_47_921 ();
 FILLCELL_X1 FILLER_47_934 ();
 FILLCELL_X4 FILLER_47_993 ();
 FILLCELL_X1 FILLER_47_997 ();
 FILLCELL_X4 FILLER_47_1003 ();
 FILLCELL_X16 FILLER_47_1039 ();
 FILLCELL_X2 FILLER_47_1084 ();
 FILLCELL_X2 FILLER_47_1144 ();
 FILLCELL_X1 FILLER_47_1146 ();
 FILLCELL_X2 FILLER_47_1166 ();
 FILLCELL_X2 FILLER_47_1233 ();
 FILLCELL_X2 FILLER_48_1 ();
 FILLCELL_X4 FILLER_48_11 ();
 FILLCELL_X2 FILLER_48_15 ();
 FILLCELL_X2 FILLER_48_21 ();
 FILLCELL_X4 FILLER_48_43 ();
 FILLCELL_X2 FILLER_48_47 ();
 FILLCELL_X1 FILLER_48_49 ();
 FILLCELL_X4 FILLER_48_70 ();
 FILLCELL_X1 FILLER_48_74 ();
 FILLCELL_X2 FILLER_48_89 ();
 FILLCELL_X1 FILLER_48_91 ();
 FILLCELL_X16 FILLER_48_106 ();
 FILLCELL_X8 FILLER_48_122 ();
 FILLCELL_X4 FILLER_48_171 ();
 FILLCELL_X1 FILLER_48_254 ();
 FILLCELL_X2 FILLER_48_322 ();
 FILLCELL_X4 FILLER_48_329 ();
 FILLCELL_X1 FILLER_48_333 ();
 FILLCELL_X8 FILLER_48_337 ();
 FILLCELL_X1 FILLER_48_352 ();
 FILLCELL_X4 FILLER_48_360 ();
 FILLCELL_X2 FILLER_48_364 ();
 FILLCELL_X1 FILLER_48_366 ();
 FILLCELL_X1 FILLER_48_380 ();
 FILLCELL_X1 FILLER_48_391 ();
 FILLCELL_X4 FILLER_48_432 ();
 FILLCELL_X2 FILLER_48_436 ();
 FILLCELL_X1 FILLER_48_438 ();
 FILLCELL_X4 FILLER_48_446 ();
 FILLCELL_X2 FILLER_48_450 ();
 FILLCELL_X1 FILLER_48_460 ();
 FILLCELL_X2 FILLER_48_470 ();
 FILLCELL_X8 FILLER_48_501 ();
 FILLCELL_X2 FILLER_48_509 ();
 FILLCELL_X4 FILLER_48_525 ();
 FILLCELL_X8 FILLER_48_549 ();
 FILLCELL_X4 FILLER_48_557 ();
 FILLCELL_X1 FILLER_48_561 ();
 FILLCELL_X1 FILLER_48_565 ();
 FILLCELL_X2 FILLER_48_573 ();
 FILLCELL_X1 FILLER_48_575 ();
 FILLCELL_X4 FILLER_48_578 ();
 FILLCELL_X2 FILLER_48_587 ();
 FILLCELL_X2 FILLER_48_596 ();
 FILLCELL_X8 FILLER_48_605 ();
 FILLCELL_X4 FILLER_48_613 ();
 FILLCELL_X2 FILLER_48_617 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X4 FILLER_48_632 ();
 FILLCELL_X1 FILLER_48_636 ();
 FILLCELL_X1 FILLER_48_646 ();
 FILLCELL_X1 FILLER_48_656 ();
 FILLCELL_X1 FILLER_48_660 ();
 FILLCELL_X4 FILLER_48_675 ();
 FILLCELL_X2 FILLER_48_679 ();
 FILLCELL_X16 FILLER_48_695 ();
 FILLCELL_X8 FILLER_48_711 ();
 FILLCELL_X16 FILLER_48_745 ();
 FILLCELL_X4 FILLER_48_780 ();
 FILLCELL_X2 FILLER_48_797 ();
 FILLCELL_X1 FILLER_48_803 ();
 FILLCELL_X2 FILLER_48_808 ();
 FILLCELL_X1 FILLER_48_810 ();
 FILLCELL_X8 FILLER_48_827 ();
 FILLCELL_X4 FILLER_48_835 ();
 FILLCELL_X1 FILLER_48_839 ();
 FILLCELL_X2 FILLER_48_846 ();
 FILLCELL_X2 FILLER_48_863 ();
 FILLCELL_X1 FILLER_48_865 ();
 FILLCELL_X2 FILLER_48_884 ();
 FILLCELL_X1 FILLER_48_886 ();
 FILLCELL_X4 FILLER_48_894 ();
 FILLCELL_X1 FILLER_48_898 ();
 FILLCELL_X8 FILLER_48_906 ();
 FILLCELL_X1 FILLER_48_914 ();
 FILLCELL_X2 FILLER_48_963 ();
 FILLCELL_X16 FILLER_48_967 ();
 FILLCELL_X8 FILLER_48_983 ();
 FILLCELL_X4 FILLER_48_991 ();
 FILLCELL_X1 FILLER_48_1008 ();
 FILLCELL_X1 FILLER_48_1022 ();
 FILLCELL_X1 FILLER_48_1026 ();
 FILLCELL_X1 FILLER_48_1031 ();
 FILLCELL_X8 FILLER_48_1035 ();
 FILLCELL_X4 FILLER_48_1043 ();
 FILLCELL_X1 FILLER_48_1047 ();
 FILLCELL_X4 FILLER_48_1068 ();
 FILLCELL_X4 FILLER_48_1119 ();
 FILLCELL_X4 FILLER_48_1134 ();
 FILLCELL_X2 FILLER_48_1138 ();
 FILLCELL_X1 FILLER_48_1140 ();
 FILLCELL_X2 FILLER_48_1148 ();
 FILLCELL_X2 FILLER_48_1188 ();
 FILLCELL_X1 FILLER_48_1190 ();
 FILLCELL_X1 FILLER_48_1195 ();
 FILLCELL_X2 FILLER_48_1199 ();
 FILLCELL_X2 FILLER_48_1208 ();
 FILLCELL_X2 FILLER_48_1226 ();
 FILLCELL_X2 FILLER_48_1253 ();
 FILLCELL_X16 FILLER_49_1 ();
 FILLCELL_X2 FILLER_49_17 ();
 FILLCELL_X1 FILLER_49_19 ();
 FILLCELL_X16 FILLER_49_28 ();
 FILLCELL_X8 FILLER_49_44 ();
 FILLCELL_X4 FILLER_49_52 ();
 FILLCELL_X1 FILLER_49_56 ();
 FILLCELL_X4 FILLER_49_64 ();
 FILLCELL_X4 FILLER_49_75 ();
 FILLCELL_X2 FILLER_49_86 ();
 FILLCELL_X1 FILLER_49_88 ();
 FILLCELL_X2 FILLER_49_117 ();
 FILLCELL_X1 FILLER_49_128 ();
 FILLCELL_X4 FILLER_49_137 ();
 FILLCELL_X2 FILLER_49_173 ();
 FILLCELL_X1 FILLER_49_175 ();
 FILLCELL_X1 FILLER_49_270 ();
 FILLCELL_X1 FILLER_49_313 ();
 FILLCELL_X2 FILLER_49_317 ();
 FILLCELL_X4 FILLER_49_344 ();
 FILLCELL_X2 FILLER_49_355 ();
 FILLCELL_X2 FILLER_49_362 ();
 FILLCELL_X4 FILLER_49_389 ();
 FILLCELL_X1 FILLER_49_393 ();
 FILLCELL_X4 FILLER_49_414 ();
 FILLCELL_X2 FILLER_49_418 ();
 FILLCELL_X1 FILLER_49_420 ();
 FILLCELL_X1 FILLER_49_446 ();
 FILLCELL_X1 FILLER_49_454 ();
 FILLCELL_X1 FILLER_49_462 ();
 FILLCELL_X1 FILLER_49_470 ();
 FILLCELL_X1 FILLER_49_478 ();
 FILLCELL_X2 FILLER_49_486 ();
 FILLCELL_X2 FILLER_49_509 ();
 FILLCELL_X1 FILLER_49_511 ();
 FILLCELL_X4 FILLER_49_533 ();
 FILLCELL_X4 FILLER_49_551 ();
 FILLCELL_X2 FILLER_49_555 ();
 FILLCELL_X1 FILLER_49_557 ();
 FILLCELL_X1 FILLER_49_592 ();
 FILLCELL_X4 FILLER_49_615 ();
 FILLCELL_X1 FILLER_49_619 ();
 FILLCELL_X2 FILLER_49_624 ();
 FILLCELL_X1 FILLER_49_626 ();
 FILLCELL_X2 FILLER_49_643 ();
 FILLCELL_X1 FILLER_49_645 ();
 FILLCELL_X1 FILLER_49_662 ();
 FILLCELL_X4 FILLER_49_681 ();
 FILLCELL_X1 FILLER_49_685 ();
 FILLCELL_X2 FILLER_49_700 ();
 FILLCELL_X8 FILLER_49_707 ();
 FILLCELL_X4 FILLER_49_715 ();
 FILLCELL_X2 FILLER_49_719 ();
 FILLCELL_X8 FILLER_49_730 ();
 FILLCELL_X2 FILLER_49_738 ();
 FILLCELL_X16 FILLER_49_769 ();
 FILLCELL_X4 FILLER_49_785 ();
 FILLCELL_X4 FILLER_49_796 ();
 FILLCELL_X1 FILLER_49_800 ();
 FILLCELL_X1 FILLER_49_809 ();
 FILLCELL_X1 FILLER_49_813 ();
 FILLCELL_X1 FILLER_49_818 ();
 FILLCELL_X1 FILLER_49_826 ();
 FILLCELL_X4 FILLER_49_844 ();
 FILLCELL_X8 FILLER_49_853 ();
 FILLCELL_X8 FILLER_49_901 ();
 FILLCELL_X4 FILLER_49_909 ();
 FILLCELL_X2 FILLER_49_913 ();
 FILLCELL_X2 FILLER_49_937 ();
 FILLCELL_X1 FILLER_49_945 ();
 FILLCELL_X4 FILLER_49_965 ();
 FILLCELL_X1 FILLER_49_969 ();
 FILLCELL_X2 FILLER_49_1022 ();
 FILLCELL_X4 FILLER_49_1067 ();
 FILLCELL_X2 FILLER_49_1078 ();
 FILLCELL_X1 FILLER_49_1091 ();
 FILLCELL_X32 FILLER_49_1110 ();
 FILLCELL_X4 FILLER_49_1142 ();
 FILLCELL_X2 FILLER_49_1146 ();
 FILLCELL_X4 FILLER_49_1162 ();
 FILLCELL_X2 FILLER_49_1166 ();
 FILLCELL_X4 FILLER_49_1182 ();
 FILLCELL_X2 FILLER_49_1186 ();
 FILLCELL_X1 FILLER_49_1195 ();
 FILLCELL_X2 FILLER_49_1219 ();
 FILLCELL_X1 FILLER_49_1221 ();
 FILLCELL_X1 FILLER_49_1250 ();
 FILLCELL_X4 FILLER_50_1 ();
 FILLCELL_X2 FILLER_50_5 ();
 FILLCELL_X2 FILLER_50_11 ();
 FILLCELL_X1 FILLER_50_13 ();
 FILLCELL_X8 FILLER_50_18 ();
 FILLCELL_X4 FILLER_50_26 ();
 FILLCELL_X2 FILLER_50_30 ();
 FILLCELL_X8 FILLER_50_40 ();
 FILLCELL_X4 FILLER_50_48 ();
 FILLCELL_X4 FILLER_50_86 ();
 FILLCELL_X1 FILLER_50_90 ();
 FILLCELL_X16 FILLER_50_98 ();
 FILLCELL_X2 FILLER_50_114 ();
 FILLCELL_X4 FILLER_50_143 ();
 FILLCELL_X1 FILLER_50_174 ();
 FILLCELL_X1 FILLER_50_326 ();
 FILLCELL_X1 FILLER_50_336 ();
 FILLCELL_X2 FILLER_50_351 ();
 FILLCELL_X2 FILLER_50_360 ();
 FILLCELL_X1 FILLER_50_362 ();
 FILLCELL_X1 FILLER_50_388 ();
 FILLCELL_X16 FILLER_50_396 ();
 FILLCELL_X8 FILLER_50_412 ();
 FILLCELL_X4 FILLER_50_420 ();
 FILLCELL_X16 FILLER_50_431 ();
 FILLCELL_X2 FILLER_50_447 ();
 FILLCELL_X2 FILLER_50_456 ();
 FILLCELL_X1 FILLER_50_470 ();
 FILLCELL_X8 FILLER_50_491 ();
 FILLCELL_X4 FILLER_50_511 ();
 FILLCELL_X1 FILLER_50_519 ();
 FILLCELL_X1 FILLER_50_559 ();
 FILLCELL_X8 FILLER_50_563 ();
 FILLCELL_X4 FILLER_50_571 ();
 FILLCELL_X1 FILLER_50_575 ();
 FILLCELL_X1 FILLER_50_583 ();
 FILLCELL_X4 FILLER_50_588 ();
 FILLCELL_X2 FILLER_50_592 ();
 FILLCELL_X2 FILLER_50_616 ();
 FILLCELL_X2 FILLER_50_628 ();
 FILLCELL_X1 FILLER_50_630 ();
 FILLCELL_X2 FILLER_50_639 ();
 FILLCELL_X2 FILLER_50_672 ();
 FILLCELL_X1 FILLER_50_686 ();
 FILLCELL_X2 FILLER_50_705 ();
 FILLCELL_X1 FILLER_50_707 ();
 FILLCELL_X4 FILLER_50_721 ();
 FILLCELL_X2 FILLER_50_725 ();
 FILLCELL_X1 FILLER_50_727 ();
 FILLCELL_X16 FILLER_50_741 ();
 FILLCELL_X1 FILLER_50_757 ();
 FILLCELL_X8 FILLER_50_763 ();
 FILLCELL_X2 FILLER_50_771 ();
 FILLCELL_X1 FILLER_50_773 ();
 FILLCELL_X2 FILLER_50_777 ();
 FILLCELL_X2 FILLER_50_788 ();
 FILLCELL_X1 FILLER_50_790 ();
 FILLCELL_X2 FILLER_50_804 ();
 FILLCELL_X1 FILLER_50_806 ();
 FILLCELL_X4 FILLER_50_810 ();
 FILLCELL_X8 FILLER_50_821 ();
 FILLCELL_X4 FILLER_50_829 ();
 FILLCELL_X1 FILLER_50_833 ();
 FILLCELL_X2 FILLER_50_837 ();
 FILLCELL_X2 FILLER_50_846 ();
 FILLCELL_X1 FILLER_50_848 ();
 FILLCELL_X1 FILLER_50_854 ();
 FILLCELL_X8 FILLER_50_872 ();
 FILLCELL_X4 FILLER_50_880 ();
 FILLCELL_X4 FILLER_50_897 ();
 FILLCELL_X8 FILLER_50_924 ();
 FILLCELL_X2 FILLER_50_932 ();
 FILLCELL_X16 FILLER_50_938 ();
 FILLCELL_X2 FILLER_50_979 ();
 FILLCELL_X8 FILLER_50_992 ();
 FILLCELL_X4 FILLER_50_1000 ();
 FILLCELL_X2 FILLER_50_1004 ();
 FILLCELL_X1 FILLER_50_1006 ();
 FILLCELL_X8 FILLER_50_1014 ();
 FILLCELL_X1 FILLER_50_1022 ();
 FILLCELL_X8 FILLER_50_1033 ();
 FILLCELL_X2 FILLER_50_1041 ();
 FILLCELL_X1 FILLER_50_1046 ();
 FILLCELL_X2 FILLER_50_1052 ();
 FILLCELL_X1 FILLER_50_1074 ();
 FILLCELL_X4 FILLER_50_1086 ();
 FILLCELL_X2 FILLER_50_1090 ();
 FILLCELL_X1 FILLER_50_1092 ();
 FILLCELL_X1 FILLER_50_1109 ();
 FILLCELL_X4 FILLER_50_1117 ();
 FILLCELL_X2 FILLER_50_1138 ();
 FILLCELL_X2 FILLER_50_1160 ();
 FILLCELL_X1 FILLER_50_1162 ();
 FILLCELL_X4 FILLER_50_1183 ();
 FILLCELL_X2 FILLER_50_1187 ();
 FILLCELL_X4 FILLER_50_1193 ();
 FILLCELL_X2 FILLER_50_1197 ();
 FILLCELL_X4 FILLER_50_1206 ();
 FILLCELL_X8 FILLER_50_1214 ();
 FILLCELL_X1 FILLER_50_1222 ();
 FILLCELL_X4 FILLER_51_1 ();
 FILLCELL_X2 FILLER_51_5 ();
 FILLCELL_X1 FILLER_51_7 ();
 FILLCELL_X2 FILLER_51_35 ();
 FILLCELL_X4 FILLER_51_75 ();
 FILLCELL_X1 FILLER_51_79 ();
 FILLCELL_X4 FILLER_51_87 ();
 FILLCELL_X1 FILLER_51_91 ();
 FILLCELL_X4 FILLER_51_108 ();
 FILLCELL_X1 FILLER_51_112 ();
 FILLCELL_X4 FILLER_51_120 ();
 FILLCELL_X2 FILLER_51_124 ();
 FILLCELL_X2 FILLER_51_164 ();
 FILLCELL_X2 FILLER_51_205 ();
 FILLCELL_X4 FILLER_51_275 ();
 FILLCELL_X2 FILLER_51_279 ();
 FILLCELL_X2 FILLER_51_317 ();
 FILLCELL_X1 FILLER_51_339 ();
 FILLCELL_X2 FILLER_51_347 ();
 FILLCELL_X4 FILLER_51_354 ();
 FILLCELL_X16 FILLER_51_361 ();
 FILLCELL_X8 FILLER_51_377 ();
 FILLCELL_X2 FILLER_51_413 ();
 FILLCELL_X1 FILLER_51_449 ();
 FILLCELL_X4 FILLER_51_509 ();
 FILLCELL_X2 FILLER_51_513 ();
 FILLCELL_X1 FILLER_51_515 ();
 FILLCELL_X8 FILLER_51_543 ();
 FILLCELL_X2 FILLER_51_551 ();
 FILLCELL_X2 FILLER_51_576 ();
 FILLCELL_X1 FILLER_51_578 ();
 FILLCELL_X4 FILLER_51_582 ();
 FILLCELL_X2 FILLER_51_586 ();
 FILLCELL_X2 FILLER_51_609 ();
 FILLCELL_X2 FILLER_51_618 ();
 FILLCELL_X2 FILLER_51_631 ();
 FILLCELL_X1 FILLER_51_633 ();
 FILLCELL_X1 FILLER_51_641 ();
 FILLCELL_X1 FILLER_51_645 ();
 FILLCELL_X1 FILLER_51_651 ();
 FILLCELL_X1 FILLER_51_659 ();
 FILLCELL_X4 FILLER_51_683 ();
 FILLCELL_X2 FILLER_51_687 ();
 FILLCELL_X1 FILLER_51_689 ();
 FILLCELL_X2 FILLER_51_709 ();
 FILLCELL_X2 FILLER_51_714 ();
 FILLCELL_X4 FILLER_51_730 ();
 FILLCELL_X4 FILLER_51_748 ();
 FILLCELL_X4 FILLER_51_776 ();
 FILLCELL_X8 FILLER_51_783 ();
 FILLCELL_X1 FILLER_51_791 ();
 FILLCELL_X16 FILLER_51_826 ();
 FILLCELL_X1 FILLER_51_842 ();
 FILLCELL_X8 FILLER_51_855 ();
 FILLCELL_X2 FILLER_51_863 ();
 FILLCELL_X1 FILLER_51_865 ();
 FILLCELL_X1 FILLER_51_882 ();
 FILLCELL_X32 FILLER_51_895 ();
 FILLCELL_X8 FILLER_51_927 ();
 FILLCELL_X4 FILLER_51_965 ();
 FILLCELL_X1 FILLER_51_969 ();
 FILLCELL_X4 FILLER_51_973 ();
 FILLCELL_X1 FILLER_51_977 ();
 FILLCELL_X8 FILLER_51_1004 ();
 FILLCELL_X1 FILLER_51_1012 ();
 FILLCELL_X2 FILLER_51_1086 ();
 FILLCELL_X8 FILLER_51_1116 ();
 FILLCELL_X2 FILLER_51_1124 ();
 FILLCELL_X8 FILLER_51_1133 ();
 FILLCELL_X2 FILLER_51_1141 ();
 FILLCELL_X4 FILLER_51_1150 ();
 FILLCELL_X2 FILLER_51_1154 ();
 FILLCELL_X1 FILLER_51_1156 ();
 FILLCELL_X2 FILLER_51_1166 ();
 FILLCELL_X16 FILLER_51_1173 ();
 FILLCELL_X4 FILLER_51_1189 ();
 FILLCELL_X2 FILLER_51_1193 ();
 FILLCELL_X1 FILLER_51_1195 ();
 FILLCELL_X2 FILLER_51_1203 ();
 FILLCELL_X1 FILLER_51_1205 ();
 FILLCELL_X1 FILLER_51_1216 ();
 FILLCELL_X1 FILLER_51_1221 ();
 FILLCELL_X8 FILLER_51_1225 ();
 FILLCELL_X1 FILLER_51_1233 ();
 FILLCELL_X1 FILLER_51_1237 ();
 FILLCELL_X2 FILLER_51_1246 ();
 FILLCELL_X1 FILLER_51_1248 ();
 FILLCELL_X2 FILLER_52_1 ();
 FILLCELL_X1 FILLER_52_3 ();
 FILLCELL_X1 FILLER_52_65 ();
 FILLCELL_X4 FILLER_52_107 ();
 FILLCELL_X1 FILLER_52_111 ();
 FILLCELL_X2 FILLER_52_132 ();
 FILLCELL_X4 FILLER_52_154 ();
 FILLCELL_X2 FILLER_52_201 ();
 FILLCELL_X4 FILLER_52_279 ();
 FILLCELL_X1 FILLER_52_290 ();
 FILLCELL_X8 FILLER_52_321 ();
 FILLCELL_X4 FILLER_52_329 ();
 FILLCELL_X1 FILLER_52_333 ();
 FILLCELL_X4 FILLER_52_381 ();
 FILLCELL_X2 FILLER_52_385 ();
 FILLCELL_X1 FILLER_52_411 ();
 FILLCELL_X4 FILLER_52_432 ();
 FILLCELL_X2 FILLER_52_436 ();
 FILLCELL_X8 FILLER_52_458 ();
 FILLCELL_X2 FILLER_52_466 ();
 FILLCELL_X1 FILLER_52_468 ();
 FILLCELL_X4 FILLER_52_483 ();
 FILLCELL_X1 FILLER_52_500 ();
 FILLCELL_X1 FILLER_52_511 ();
 FILLCELL_X2 FILLER_52_534 ();
 FILLCELL_X1 FILLER_52_536 ();
 FILLCELL_X1 FILLER_52_550 ();
 FILLCELL_X2 FILLER_52_570 ();
 FILLCELL_X1 FILLER_52_587 ();
 FILLCELL_X2 FILLER_52_591 ();
 FILLCELL_X16 FILLER_52_602 ();
 FILLCELL_X8 FILLER_52_618 ();
 FILLCELL_X4 FILLER_52_626 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X4 FILLER_52_657 ();
 FILLCELL_X1 FILLER_52_661 ();
 FILLCELL_X8 FILLER_52_671 ();
 FILLCELL_X1 FILLER_52_716 ();
 FILLCELL_X8 FILLER_52_721 ();
 FILLCELL_X2 FILLER_52_729 ();
 FILLCELL_X8 FILLER_52_738 ();
 FILLCELL_X4 FILLER_52_746 ();
 FILLCELL_X4 FILLER_52_768 ();
 FILLCELL_X1 FILLER_52_797 ();
 FILLCELL_X2 FILLER_52_812 ();
 FILLCELL_X4 FILLER_52_828 ();
 FILLCELL_X2 FILLER_52_832 ();
 FILLCELL_X8 FILLER_52_857 ();
 FILLCELL_X2 FILLER_52_865 ();
 FILLCELL_X1 FILLER_52_867 ();
 FILLCELL_X4 FILLER_52_875 ();
 FILLCELL_X2 FILLER_52_879 ();
 FILLCELL_X4 FILLER_52_894 ();
 FILLCELL_X1 FILLER_52_918 ();
 FILLCELL_X1 FILLER_52_922 ();
 FILLCELL_X1 FILLER_52_930 ();
 FILLCELL_X1 FILLER_52_936 ();
 FILLCELL_X2 FILLER_52_947 ();
 FILLCELL_X4 FILLER_52_956 ();
 FILLCELL_X4 FILLER_52_962 ();
 FILLCELL_X2 FILLER_52_966 ();
 FILLCELL_X1 FILLER_52_968 ();
 FILLCELL_X8 FILLER_52_976 ();
 FILLCELL_X4 FILLER_52_984 ();
 FILLCELL_X2 FILLER_52_988 ();
 FILLCELL_X1 FILLER_52_990 ();
 FILLCELL_X8 FILLER_52_1016 ();
 FILLCELL_X2 FILLER_52_1024 ();
 FILLCELL_X1 FILLER_52_1026 ();
 FILLCELL_X8 FILLER_52_1033 ();
 FILLCELL_X4 FILLER_52_1041 ();
 FILLCELL_X1 FILLER_52_1045 ();
 FILLCELL_X1 FILLER_52_1049 ();
 FILLCELL_X2 FILLER_52_1055 ();
 FILLCELL_X16 FILLER_52_1065 ();
 FILLCELL_X4 FILLER_52_1081 ();
 FILLCELL_X2 FILLER_52_1085 ();
 FILLCELL_X1 FILLER_52_1087 ();
 FILLCELL_X2 FILLER_52_1118 ();
 FILLCELL_X4 FILLER_52_1149 ();
 FILLCELL_X8 FILLER_52_1162 ();
 FILLCELL_X4 FILLER_52_1170 ();
 FILLCELL_X2 FILLER_52_1174 ();
 FILLCELL_X1 FILLER_52_1176 ();
 FILLCELL_X2 FILLER_52_1195 ();
 FILLCELL_X4 FILLER_52_1227 ();
 FILLCELL_X1 FILLER_52_1231 ();
 FILLCELL_X1 FILLER_52_1254 ();
 FILLCELL_X8 FILLER_53_1 ();
 FILLCELL_X4 FILLER_53_9 ();
 FILLCELL_X2 FILLER_53_13 ();
 FILLCELL_X16 FILLER_53_22 ();
 FILLCELL_X8 FILLER_53_38 ();
 FILLCELL_X4 FILLER_53_46 ();
 FILLCELL_X2 FILLER_53_90 ();
 FILLCELL_X1 FILLER_53_92 ();
 FILLCELL_X4 FILLER_53_141 ();
 FILLCELL_X2 FILLER_53_145 ();
 FILLCELL_X1 FILLER_53_174 ();
 FILLCELL_X2 FILLER_53_236 ();
 FILLCELL_X2 FILLER_53_278 ();
 FILLCELL_X1 FILLER_53_287 ();
 FILLCELL_X2 FILLER_53_295 ();
 FILLCELL_X2 FILLER_53_304 ();
 FILLCELL_X1 FILLER_53_306 ();
 FILLCELL_X1 FILLER_53_331 ();
 FILLCELL_X2 FILLER_53_388 ();
 FILLCELL_X4 FILLER_53_400 ();
 FILLCELL_X2 FILLER_53_404 ();
 FILLCELL_X8 FILLER_53_420 ();
 FILLCELL_X2 FILLER_53_428 ();
 FILLCELL_X1 FILLER_53_430 ();
 FILLCELL_X1 FILLER_53_479 ();
 FILLCELL_X4 FILLER_53_482 ();
 FILLCELL_X4 FILLER_53_490 ();
 FILLCELL_X32 FILLER_53_510 ();
 FILLCELL_X8 FILLER_53_542 ();
 FILLCELL_X4 FILLER_53_550 ();
 FILLCELL_X1 FILLER_53_554 ();
 FILLCELL_X1 FILLER_53_557 ();
 FILLCELL_X4 FILLER_53_569 ();
 FILLCELL_X4 FILLER_53_576 ();
 FILLCELL_X1 FILLER_53_580 ();
 FILLCELL_X1 FILLER_53_591 ();
 FILLCELL_X16 FILLER_53_600 ();
 FILLCELL_X4 FILLER_53_616 ();
 FILLCELL_X2 FILLER_53_634 ();
 FILLCELL_X1 FILLER_53_636 ();
 FILLCELL_X2 FILLER_53_646 ();
 FILLCELL_X1 FILLER_53_648 ();
 FILLCELL_X1 FILLER_53_675 ();
 FILLCELL_X4 FILLER_53_692 ();
 FILLCELL_X2 FILLER_53_696 ();
 FILLCELL_X1 FILLER_53_698 ();
 FILLCELL_X1 FILLER_53_710 ();
 FILLCELL_X2 FILLER_53_723 ();
 FILLCELL_X2 FILLER_53_730 ();
 FILLCELL_X1 FILLER_53_732 ();
 FILLCELL_X2 FILLER_53_753 ();
 FILLCELL_X1 FILLER_53_755 ();
 FILLCELL_X2 FILLER_53_760 ();
 FILLCELL_X1 FILLER_53_765 ();
 FILLCELL_X1 FILLER_53_773 ();
 FILLCELL_X2 FILLER_53_778 ();
 FILLCELL_X4 FILLER_53_792 ();
 FILLCELL_X1 FILLER_53_796 ();
 FILLCELL_X4 FILLER_53_812 ();
 FILLCELL_X8 FILLER_53_833 ();
 FILLCELL_X2 FILLER_53_841 ();
 FILLCELL_X1 FILLER_53_843 ();
 FILLCELL_X2 FILLER_53_873 ();
 FILLCELL_X1 FILLER_53_875 ();
 FILLCELL_X2 FILLER_53_883 ();
 FILLCELL_X1 FILLER_53_885 ();
 FILLCELL_X2 FILLER_53_893 ();
 FILLCELL_X2 FILLER_53_902 ();
 FILLCELL_X1 FILLER_53_904 ();
 FILLCELL_X1 FILLER_53_909 ();
 FILLCELL_X2 FILLER_53_917 ();
 FILLCELL_X1 FILLER_53_919 ();
 FILLCELL_X1 FILLER_53_924 ();
 FILLCELL_X16 FILLER_53_936 ();
 FILLCELL_X1 FILLER_53_952 ();
 FILLCELL_X2 FILLER_53_956 ();
 FILLCELL_X1 FILLER_53_958 ();
 FILLCELL_X2 FILLER_53_969 ();
 FILLCELL_X2 FILLER_53_994 ();
 FILLCELL_X1 FILLER_53_1016 ();
 FILLCELL_X4 FILLER_53_1037 ();
 FILLCELL_X2 FILLER_53_1041 ();
 FILLCELL_X1 FILLER_53_1043 ();
 FILLCELL_X1 FILLER_53_1051 ();
 FILLCELL_X1 FILLER_53_1054 ();
 FILLCELL_X4 FILLER_53_1063 ();
 FILLCELL_X1 FILLER_53_1067 ();
 FILLCELL_X1 FILLER_53_1077 ();
 FILLCELL_X2 FILLER_53_1098 ();
 FILLCELL_X1 FILLER_53_1100 ();
 FILLCELL_X16 FILLER_53_1119 ();
 FILLCELL_X1 FILLER_53_1135 ();
 FILLCELL_X1 FILLER_53_1156 ();
 FILLCELL_X4 FILLER_53_1179 ();
 FILLCELL_X1 FILLER_53_1183 ();
 FILLCELL_X2 FILLER_53_1208 ();
 FILLCELL_X1 FILLER_53_1210 ();
 FILLCELL_X4 FILLER_53_1218 ();
 FILLCELL_X2 FILLER_53_1253 ();
 FILLCELL_X16 FILLER_54_48 ();
 FILLCELL_X8 FILLER_54_64 ();
 FILLCELL_X4 FILLER_54_72 ();
 FILLCELL_X4 FILLER_54_90 ();
 FILLCELL_X2 FILLER_54_94 ();
 FILLCELL_X2 FILLER_54_110 ();
 FILLCELL_X2 FILLER_54_119 ();
 FILLCELL_X16 FILLER_54_135 ();
 FILLCELL_X1 FILLER_54_286 ();
 FILLCELL_X2 FILLER_54_310 ();
 FILLCELL_X1 FILLER_54_318 ();
 FILLCELL_X2 FILLER_54_329 ();
 FILLCELL_X1 FILLER_54_331 ();
 FILLCELL_X4 FILLER_54_346 ();
 FILLCELL_X2 FILLER_54_350 ();
 FILLCELL_X2 FILLER_54_368 ();
 FILLCELL_X2 FILLER_54_380 ();
 FILLCELL_X1 FILLER_54_382 ();
 FILLCELL_X2 FILLER_54_417 ();
 FILLCELL_X4 FILLER_54_426 ();
 FILLCELL_X2 FILLER_54_430 ();
 FILLCELL_X1 FILLER_54_432 ();
 FILLCELL_X4 FILLER_54_466 ();
 FILLCELL_X2 FILLER_54_470 ();
 FILLCELL_X4 FILLER_54_487 ();
 FILLCELL_X2 FILLER_54_498 ();
 FILLCELL_X1 FILLER_54_500 ();
 FILLCELL_X8 FILLER_54_503 ();
 FILLCELL_X4 FILLER_54_511 ();
 FILLCELL_X8 FILLER_54_520 ();
 FILLCELL_X1 FILLER_54_553 ();
 FILLCELL_X2 FILLER_54_568 ();
 FILLCELL_X1 FILLER_54_570 ();
 FILLCELL_X1 FILLER_54_607 ();
 FILLCELL_X8 FILLER_54_610 ();
 FILLCELL_X8 FILLER_54_623 ();
 FILLCELL_X2 FILLER_54_632 ();
 FILLCELL_X4 FILLER_54_647 ();
 FILLCELL_X4 FILLER_54_658 ();
 FILLCELL_X2 FILLER_54_673 ();
 FILLCELL_X1 FILLER_54_675 ();
 FILLCELL_X2 FILLER_54_692 ();
 FILLCELL_X1 FILLER_54_698 ();
 FILLCELL_X2 FILLER_54_728 ();
 FILLCELL_X1 FILLER_54_730 ();
 FILLCELL_X4 FILLER_54_736 ();
 FILLCELL_X2 FILLER_54_740 ();
 FILLCELL_X2 FILLER_54_753 ();
 FILLCELL_X1 FILLER_54_755 ();
 FILLCELL_X1 FILLER_54_761 ();
 FILLCELL_X2 FILLER_54_769 ();
 FILLCELL_X1 FILLER_54_771 ();
 FILLCELL_X4 FILLER_54_784 ();
 FILLCELL_X1 FILLER_54_790 ();
 FILLCELL_X16 FILLER_54_819 ();
 FILLCELL_X4 FILLER_54_835 ();
 FILLCELL_X16 FILLER_54_853 ();
 FILLCELL_X4 FILLER_54_869 ();
 FILLCELL_X16 FILLER_54_912 ();
 FILLCELL_X1 FILLER_54_928 ();
 FILLCELL_X8 FILLER_54_938 ();
 FILLCELL_X1 FILLER_54_946 ();
 FILLCELL_X1 FILLER_54_961 ();
 FILLCELL_X2 FILLER_54_967 ();
 FILLCELL_X1 FILLER_54_969 ();
 FILLCELL_X2 FILLER_54_997 ();
 FILLCELL_X1 FILLER_54_999 ();
 FILLCELL_X1 FILLER_54_1012 ();
 FILLCELL_X8 FILLER_54_1022 ();
 FILLCELL_X2 FILLER_54_1030 ();
 FILLCELL_X1 FILLER_54_1032 ();
 FILLCELL_X1 FILLER_54_1077 ();
 FILLCELL_X8 FILLER_54_1141 ();
 FILLCELL_X4 FILLER_54_1149 ();
 FILLCELL_X1 FILLER_54_1153 ();
 FILLCELL_X4 FILLER_54_1162 ();
 FILLCELL_X2 FILLER_54_1175 ();
 FILLCELL_X8 FILLER_54_1184 ();
 FILLCELL_X1 FILLER_54_1192 ();
 FILLCELL_X4 FILLER_54_1196 ();
 FILLCELL_X1 FILLER_54_1200 ();
 FILLCELL_X2 FILLER_54_1213 ();
 FILLCELL_X1 FILLER_54_1215 ();
 FILLCELL_X1 FILLER_54_1224 ();
 FILLCELL_X4 FILLER_54_1228 ();
 FILLCELL_X1 FILLER_54_1232 ();
 FILLCELL_X2 FILLER_54_1253 ();
 FILLCELL_X4 FILLER_55_9 ();
 FILLCELL_X1 FILLER_55_13 ();
 FILLCELL_X2 FILLER_55_21 ();
 FILLCELL_X1 FILLER_55_23 ();
 FILLCELL_X8 FILLER_55_51 ();
 FILLCELL_X1 FILLER_55_71 ();
 FILLCELL_X4 FILLER_55_119 ();
 FILLCELL_X4 FILLER_55_130 ();
 FILLCELL_X1 FILLER_55_148 ();
 FILLCELL_X2 FILLER_55_169 ();
 FILLCELL_X8 FILLER_55_346 ();
 FILLCELL_X2 FILLER_55_374 ();
 FILLCELL_X2 FILLER_55_383 ();
 FILLCELL_X1 FILLER_55_385 ();
 FILLCELL_X4 FILLER_55_393 ();
 FILLCELL_X2 FILLER_55_397 ();
 FILLCELL_X1 FILLER_55_399 ();
 FILLCELL_X2 FILLER_55_421 ();
 FILLCELL_X1 FILLER_55_430 ();
 FILLCELL_X1 FILLER_55_442 ();
 FILLCELL_X1 FILLER_55_458 ();
 FILLCELL_X1 FILLER_55_464 ();
 FILLCELL_X8 FILLER_55_483 ();
 FILLCELL_X4 FILLER_55_491 ();
 FILLCELL_X2 FILLER_55_495 ();
 FILLCELL_X1 FILLER_55_497 ();
 FILLCELL_X8 FILLER_55_511 ();
 FILLCELL_X4 FILLER_55_519 ();
 FILLCELL_X2 FILLER_55_523 ();
 FILLCELL_X1 FILLER_55_525 ();
 FILLCELL_X1 FILLER_55_553 ();
 FILLCELL_X4 FILLER_55_562 ();
 FILLCELL_X4 FILLER_55_568 ();
 FILLCELL_X8 FILLER_55_588 ();
 FILLCELL_X1 FILLER_55_596 ();
 FILLCELL_X32 FILLER_55_604 ();
 FILLCELL_X1 FILLER_55_636 ();
 FILLCELL_X4 FILLER_55_649 ();
 FILLCELL_X1 FILLER_55_653 ();
 FILLCELL_X4 FILLER_55_689 ();
 FILLCELL_X1 FILLER_55_693 ();
 FILLCELL_X2 FILLER_55_717 ();
 FILLCELL_X1 FILLER_55_719 ();
 FILLCELL_X4 FILLER_55_724 ();
 FILLCELL_X4 FILLER_55_754 ();
 FILLCELL_X2 FILLER_55_758 ();
 FILLCELL_X1 FILLER_55_760 ();
 FILLCELL_X2 FILLER_55_770 ();
 FILLCELL_X1 FILLER_55_772 ();
 FILLCELL_X8 FILLER_55_778 ();
 FILLCELL_X1 FILLER_55_786 ();
 FILLCELL_X2 FILLER_55_791 ();
 FILLCELL_X2 FILLER_55_800 ();
 FILLCELL_X1 FILLER_55_802 ();
 FILLCELL_X4 FILLER_55_810 ();
 FILLCELL_X1 FILLER_55_814 ();
 FILLCELL_X2 FILLER_55_835 ();
 FILLCELL_X2 FILLER_55_851 ();
 FILLCELL_X4 FILLER_55_864 ();
 FILLCELL_X1 FILLER_55_868 ();
 FILLCELL_X4 FILLER_55_874 ();
 FILLCELL_X2 FILLER_55_878 ();
 FILLCELL_X2 FILLER_55_889 ();
 FILLCELL_X1 FILLER_55_927 ();
 FILLCELL_X8 FILLER_55_944 ();
 FILLCELL_X16 FILLER_55_966 ();
 FILLCELL_X4 FILLER_55_989 ();
 FILLCELL_X1 FILLER_55_993 ();
 FILLCELL_X2 FILLER_55_997 ();
 FILLCELL_X4 FILLER_55_1006 ();
 FILLCELL_X2 FILLER_55_1010 ();
 FILLCELL_X1 FILLER_55_1012 ();
 FILLCELL_X8 FILLER_55_1019 ();
 FILLCELL_X2 FILLER_55_1027 ();
 FILLCELL_X8 FILLER_55_1040 ();
 FILLCELL_X8 FILLER_55_1062 ();
 FILLCELL_X1 FILLER_55_1079 ();
 FILLCELL_X4 FILLER_55_1102 ();
 FILLCELL_X2 FILLER_55_1106 ();
 FILLCELL_X4 FILLER_55_1110 ();
 FILLCELL_X1 FILLER_55_1114 ();
 FILLCELL_X2 FILLER_55_1120 ();
 FILLCELL_X2 FILLER_55_1129 ();
 FILLCELL_X1 FILLER_55_1131 ();
 FILLCELL_X4 FILLER_55_1149 ();
 FILLCELL_X1 FILLER_55_1153 ();
 FILLCELL_X2 FILLER_55_1161 ();
 FILLCELL_X1 FILLER_55_1169 ();
 FILLCELL_X1 FILLER_55_1190 ();
 FILLCELL_X1 FILLER_55_1215 ();
 FILLCELL_X1 FILLER_55_1222 ();
 FILLCELL_X2 FILLER_55_1249 ();
 FILLCELL_X1 FILLER_55_1251 ();
 FILLCELL_X2 FILLER_56_1 ();
 FILLCELL_X1 FILLER_56_34 ();
 FILLCELL_X8 FILLER_56_39 ();
 FILLCELL_X4 FILLER_56_47 ();
 FILLCELL_X1 FILLER_56_64 ();
 FILLCELL_X1 FILLER_56_106 ();
 FILLCELL_X1 FILLER_56_119 ();
 FILLCELL_X2 FILLER_56_134 ();
 FILLCELL_X8 FILLER_56_143 ();
 FILLCELL_X1 FILLER_56_151 ();
 FILLCELL_X2 FILLER_56_247 ();
 FILLCELL_X1 FILLER_56_249 ();
 FILLCELL_X2 FILLER_56_278 ();
 FILLCELL_X1 FILLER_56_287 ();
 FILLCELL_X2 FILLER_56_293 ();
 FILLCELL_X4 FILLER_56_355 ();
 FILLCELL_X2 FILLER_56_372 ();
 FILLCELL_X1 FILLER_56_374 ();
 FILLCELL_X4 FILLER_56_396 ();
 FILLCELL_X1 FILLER_56_414 ();
 FILLCELL_X4 FILLER_56_436 ();
 FILLCELL_X2 FILLER_56_440 ();
 FILLCELL_X1 FILLER_56_442 ();
 FILLCELL_X2 FILLER_56_460 ();
 FILLCELL_X4 FILLER_56_475 ();
 FILLCELL_X1 FILLER_56_479 ();
 FILLCELL_X2 FILLER_56_487 ();
 FILLCELL_X1 FILLER_56_489 ();
 FILLCELL_X4 FILLER_56_503 ();
 FILLCELL_X1 FILLER_56_516 ();
 FILLCELL_X8 FILLER_56_543 ();
 FILLCELL_X1 FILLER_56_551 ();
 FILLCELL_X1 FILLER_56_555 ();
 FILLCELL_X4 FILLER_56_581 ();
 FILLCELL_X1 FILLER_56_585 ();
 FILLCELL_X8 FILLER_56_612 ();
 FILLCELL_X4 FILLER_56_620 ();
 FILLCELL_X1 FILLER_56_624 ();
 FILLCELL_X1 FILLER_56_630 ();
 FILLCELL_X1 FILLER_56_637 ();
 FILLCELL_X8 FILLER_56_645 ();
 FILLCELL_X2 FILLER_56_653 ();
 FILLCELL_X1 FILLER_56_672 ();
 FILLCELL_X2 FILLER_56_694 ();
 FILLCELL_X4 FILLER_56_735 ();
 FILLCELL_X2 FILLER_56_739 ();
 FILLCELL_X1 FILLER_56_741 ();
 FILLCELL_X2 FILLER_56_784 ();
 FILLCELL_X1 FILLER_56_786 ();
 FILLCELL_X2 FILLER_56_792 ();
 FILLCELL_X1 FILLER_56_794 ();
 FILLCELL_X1 FILLER_56_821 ();
 FILLCELL_X2 FILLER_56_827 ();
 FILLCELL_X1 FILLER_56_829 ();
 FILLCELL_X8 FILLER_56_834 ();
 FILLCELL_X4 FILLER_56_859 ();
 FILLCELL_X1 FILLER_56_863 ();
 FILLCELL_X4 FILLER_56_872 ();
 FILLCELL_X1 FILLER_56_876 ();
 FILLCELL_X4 FILLER_56_901 ();
 FILLCELL_X2 FILLER_56_905 ();
 FILLCELL_X4 FILLER_56_916 ();
 FILLCELL_X1 FILLER_56_920 ();
 FILLCELL_X4 FILLER_56_928 ();
 FILLCELL_X2 FILLER_56_932 ();
 FILLCELL_X4 FILLER_56_942 ();
 FILLCELL_X2 FILLER_56_951 ();
 FILLCELL_X1 FILLER_56_953 ();
 FILLCELL_X2 FILLER_56_961 ();
 FILLCELL_X4 FILLER_56_1009 ();
 FILLCELL_X1 FILLER_56_1022 ();
 FILLCELL_X2 FILLER_56_1025 ();
 FILLCELL_X4 FILLER_56_1055 ();
 FILLCELL_X2 FILLER_56_1059 ();
 FILLCELL_X1 FILLER_56_1061 ();
 FILLCELL_X2 FILLER_56_1067 ();
 FILLCELL_X1 FILLER_56_1069 ();
 FILLCELL_X1 FILLER_56_1075 ();
 FILLCELL_X2 FILLER_56_1081 ();
 FILLCELL_X1 FILLER_56_1083 ();
 FILLCELL_X4 FILLER_56_1110 ();
 FILLCELL_X2 FILLER_56_1136 ();
 FILLCELL_X4 FILLER_56_1145 ();
 FILLCELL_X4 FILLER_56_1156 ();
 FILLCELL_X1 FILLER_56_1163 ();
 FILLCELL_X1 FILLER_56_1167 ();
 FILLCELL_X2 FILLER_56_1175 ();
 FILLCELL_X4 FILLER_56_1180 ();
 FILLCELL_X2 FILLER_56_1184 ();
 FILLCELL_X2 FILLER_56_1223 ();
 FILLCELL_X1 FILLER_56_1225 ();
 FILLCELL_X2 FILLER_56_1233 ();
 FILLCELL_X4 FILLER_56_1238 ();
 FILLCELL_X2 FILLER_56_1242 ();
 FILLCELL_X2 FILLER_57_5 ();
 FILLCELL_X2 FILLER_57_36 ();
 FILLCELL_X1 FILLER_57_45 ();
 FILLCELL_X1 FILLER_57_53 ();
 FILLCELL_X1 FILLER_57_74 ();
 FILLCELL_X2 FILLER_57_82 ();
 FILLCELL_X2 FILLER_57_91 ();
 FILLCELL_X1 FILLER_57_93 ();
 FILLCELL_X1 FILLER_57_101 ();
 FILLCELL_X8 FILLER_57_143 ();
 FILLCELL_X4 FILLER_57_151 ();
 FILLCELL_X2 FILLER_57_155 ();
 FILLCELL_X1 FILLER_57_177 ();
 FILLCELL_X2 FILLER_57_262 ();
 FILLCELL_X1 FILLER_57_312 ();
 FILLCELL_X2 FILLER_57_333 ();
 FILLCELL_X1 FILLER_57_335 ();
 FILLCELL_X2 FILLER_57_350 ();
 FILLCELL_X4 FILLER_57_392 ();
 FILLCELL_X2 FILLER_57_396 ();
 FILLCELL_X8 FILLER_57_405 ();
 FILLCELL_X4 FILLER_57_425 ();
 FILLCELL_X1 FILLER_57_429 ();
 FILLCELL_X8 FILLER_57_437 ();
 FILLCELL_X4 FILLER_57_445 ();
 FILLCELL_X2 FILLER_57_449 ();
 FILLCELL_X1 FILLER_57_483 ();
 FILLCELL_X4 FILLER_57_487 ();
 FILLCELL_X2 FILLER_57_491 ();
 FILLCELL_X1 FILLER_57_493 ();
 FILLCELL_X2 FILLER_57_519 ();
 FILLCELL_X1 FILLER_57_521 ();
 FILLCELL_X4 FILLER_57_532 ();
 FILLCELL_X1 FILLER_57_536 ();
 FILLCELL_X2 FILLER_57_555 ();
 FILLCELL_X2 FILLER_57_568 ();
 FILLCELL_X1 FILLER_57_570 ();
 FILLCELL_X4 FILLER_57_595 ();
 FILLCELL_X1 FILLER_57_599 ();
 FILLCELL_X1 FILLER_57_616 ();
 FILLCELL_X4 FILLER_57_626 ();
 FILLCELL_X2 FILLER_57_630 ();
 FILLCELL_X2 FILLER_57_636 ();
 FILLCELL_X1 FILLER_57_638 ();
 FILLCELL_X1 FILLER_57_661 ();
 FILLCELL_X4 FILLER_57_683 ();
 FILLCELL_X2 FILLER_57_687 ();
 FILLCELL_X8 FILLER_57_709 ();
 FILLCELL_X2 FILLER_57_717 ();
 FILLCELL_X1 FILLER_57_722 ();
 FILLCELL_X4 FILLER_57_736 ();
 FILLCELL_X2 FILLER_57_740 ();
 FILLCELL_X1 FILLER_57_742 ();
 FILLCELL_X4 FILLER_57_746 ();
 FILLCELL_X2 FILLER_57_750 ();
 FILLCELL_X1 FILLER_57_752 ();
 FILLCELL_X8 FILLER_57_777 ();
 FILLCELL_X4 FILLER_57_802 ();
 FILLCELL_X1 FILLER_57_806 ();
 FILLCELL_X4 FILLER_57_816 ();
 FILLCELL_X1 FILLER_57_847 ();
 FILLCELL_X8 FILLER_57_852 ();
 FILLCELL_X2 FILLER_57_860 ();
 FILLCELL_X16 FILLER_57_870 ();
 FILLCELL_X8 FILLER_57_886 ();
 FILLCELL_X4 FILLER_57_894 ();
 FILLCELL_X4 FILLER_57_903 ();
 FILLCELL_X2 FILLER_57_907 ();
 FILLCELL_X1 FILLER_57_918 ();
 FILLCELL_X2 FILLER_57_927 ();
 FILLCELL_X1 FILLER_57_973 ();
 FILLCELL_X8 FILLER_57_989 ();
 FILLCELL_X1 FILLER_57_997 ();
 FILLCELL_X2 FILLER_57_1002 ();
 FILLCELL_X2 FILLER_57_1025 ();
 FILLCELL_X2 FILLER_57_1036 ();
 FILLCELL_X1 FILLER_57_1038 ();
 FILLCELL_X2 FILLER_57_1044 ();
 FILLCELL_X4 FILLER_57_1057 ();
 FILLCELL_X1 FILLER_57_1061 ();
 FILLCELL_X4 FILLER_57_1071 ();
 FILLCELL_X2 FILLER_57_1075 ();
 FILLCELL_X1 FILLER_57_1077 ();
 FILLCELL_X8 FILLER_57_1086 ();
 FILLCELL_X2 FILLER_57_1094 ();
 FILLCELL_X1 FILLER_57_1107 ();
 FILLCELL_X4 FILLER_57_1111 ();
 FILLCELL_X4 FILLER_57_1148 ();
 FILLCELL_X8 FILLER_57_1172 ();
 FILLCELL_X8 FILLER_57_1189 ();
 FILLCELL_X4 FILLER_57_1201 ();
 FILLCELL_X1 FILLER_57_1205 ();
 FILLCELL_X4 FILLER_57_1209 ();
 FILLCELL_X1 FILLER_57_1234 ();
 FILLCELL_X2 FILLER_58_1 ();
 FILLCELL_X8 FILLER_58_41 ();
 FILLCELL_X2 FILLER_58_89 ();
 FILLCELL_X2 FILLER_58_105 ();
 FILLCELL_X1 FILLER_58_177 ();
 FILLCELL_X1 FILLER_58_279 ();
 FILLCELL_X4 FILLER_58_287 ();
 FILLCELL_X2 FILLER_58_291 ();
 FILLCELL_X2 FILLER_58_325 ();
 FILLCELL_X2 FILLER_58_352 ();
 FILLCELL_X1 FILLER_58_354 ();
 FILLCELL_X2 FILLER_58_398 ();
 FILLCELL_X16 FILLER_58_403 ();
 FILLCELL_X8 FILLER_58_440 ();
 FILLCELL_X4 FILLER_58_448 ();
 FILLCELL_X16 FILLER_58_459 ();
 FILLCELL_X4 FILLER_58_475 ();
 FILLCELL_X2 FILLER_58_479 ();
 FILLCELL_X4 FILLER_58_488 ();
 FILLCELL_X8 FILLER_58_504 ();
 FILLCELL_X4 FILLER_58_512 ();
 FILLCELL_X1 FILLER_58_516 ();
 FILLCELL_X1 FILLER_58_563 ();
 FILLCELL_X1 FILLER_58_568 ();
 FILLCELL_X8 FILLER_58_571 ();
 FILLCELL_X4 FILLER_58_579 ();
 FILLCELL_X2 FILLER_58_583 ();
 FILLCELL_X1 FILLER_58_585 ();
 FILLCELL_X8 FILLER_58_592 ();
 FILLCELL_X2 FILLER_58_600 ();
 FILLCELL_X4 FILLER_58_616 ();
 FILLCELL_X4 FILLER_58_627 ();
 FILLCELL_X2 FILLER_58_643 ();
 FILLCELL_X4 FILLER_58_652 ();
 FILLCELL_X1 FILLER_58_656 ();
 FILLCELL_X4 FILLER_58_664 ();
 FILLCELL_X2 FILLER_58_668 ();
 FILLCELL_X32 FILLER_58_677 ();
 FILLCELL_X8 FILLER_58_709 ();
 FILLCELL_X2 FILLER_58_717 ();
 FILLCELL_X2 FILLER_58_762 ();
 FILLCELL_X1 FILLER_58_764 ();
 FILLCELL_X4 FILLER_58_769 ();
 FILLCELL_X2 FILLER_58_773 ();
 FILLCELL_X16 FILLER_58_781 ();
 FILLCELL_X1 FILLER_58_797 ();
 FILLCELL_X4 FILLER_58_803 ();
 FILLCELL_X1 FILLER_58_828 ();
 FILLCELL_X1 FILLER_58_833 ();
 FILLCELL_X4 FILLER_58_854 ();
 FILLCELL_X2 FILLER_58_858 ();
 FILLCELL_X8 FILLER_58_873 ();
 FILLCELL_X4 FILLER_58_881 ();
 FILLCELL_X2 FILLER_58_885 ();
 FILLCELL_X1 FILLER_58_887 ();
 FILLCELL_X8 FILLER_58_905 ();
 FILLCELL_X4 FILLER_58_913 ();
 FILLCELL_X1 FILLER_58_917 ();
 FILLCELL_X2 FILLER_58_921 ();
 FILLCELL_X4 FILLER_58_925 ();
 FILLCELL_X2 FILLER_58_929 ();
 FILLCELL_X8 FILLER_58_934 ();
 FILLCELL_X2 FILLER_58_942 ();
 FILLCELL_X8 FILLER_58_955 ();
 FILLCELL_X4 FILLER_58_967 ();
 FILLCELL_X16 FILLER_58_974 ();
 FILLCELL_X2 FILLER_58_990 ();
 FILLCELL_X2 FILLER_58_1012 ();
 FILLCELL_X2 FILLER_58_1019 ();
 FILLCELL_X2 FILLER_58_1052 ();
 FILLCELL_X1 FILLER_58_1054 ();
 FILLCELL_X2 FILLER_58_1061 ();
 FILLCELL_X1 FILLER_58_1063 ();
 FILLCELL_X4 FILLER_58_1094 ();
 FILLCELL_X2 FILLER_58_1114 ();
 FILLCELL_X1 FILLER_58_1116 ();
 FILLCELL_X8 FILLER_58_1176 ();
 FILLCELL_X4 FILLER_58_1184 ();
 FILLCELL_X2 FILLER_58_1188 ();
 FILLCELL_X1 FILLER_58_1190 ();
 FILLCELL_X8 FILLER_58_1218 ();
 FILLCELL_X2 FILLER_58_1226 ();
 FILLCELL_X1 FILLER_59_1 ();
 FILLCELL_X2 FILLER_59_29 ();
 FILLCELL_X8 FILLER_59_59 ();
 FILLCELL_X4 FILLER_59_67 ();
 FILLCELL_X1 FILLER_59_91 ();
 FILLCELL_X8 FILLER_59_99 ();
 FILLCELL_X4 FILLER_59_107 ();
 FILLCELL_X2 FILLER_59_111 ();
 FILLCELL_X1 FILLER_59_113 ();
 FILLCELL_X4 FILLER_59_121 ();
 FILLCELL_X1 FILLER_59_125 ();
 FILLCELL_X2 FILLER_59_140 ();
 FILLCELL_X1 FILLER_59_142 ();
 FILLCELL_X16 FILLER_59_157 ();
 FILLCELL_X4 FILLER_59_173 ();
 FILLCELL_X2 FILLER_59_179 ();
 FILLCELL_X1 FILLER_59_273 ();
 FILLCELL_X2 FILLER_59_301 ();
 FILLCELL_X1 FILLER_59_354 ();
 FILLCELL_X2 FILLER_59_406 ();
 FILLCELL_X4 FILLER_59_411 ();
 FILLCELL_X1 FILLER_59_415 ();
 FILLCELL_X1 FILLER_59_420 ();
 FILLCELL_X8 FILLER_59_431 ();
 FILLCELL_X2 FILLER_59_439 ();
 FILLCELL_X2 FILLER_59_455 ();
 FILLCELL_X8 FILLER_59_477 ();
 FILLCELL_X2 FILLER_59_485 ();
 FILLCELL_X1 FILLER_59_487 ();
 FILLCELL_X4 FILLER_59_500 ();
 FILLCELL_X2 FILLER_59_504 ();
 FILLCELL_X2 FILLER_59_509 ();
 FILLCELL_X1 FILLER_59_511 ();
 FILLCELL_X4 FILLER_59_539 ();
 FILLCELL_X2 FILLER_59_543 ();
 FILLCELL_X1 FILLER_59_545 ();
 FILLCELL_X1 FILLER_59_558 ();
 FILLCELL_X8 FILLER_59_570 ();
 FILLCELL_X2 FILLER_59_596 ();
 FILLCELL_X2 FILLER_59_607 ();
 FILLCELL_X8 FILLER_59_632 ();
 FILLCELL_X4 FILLER_59_640 ();
 FILLCELL_X1 FILLER_59_644 ();
 FILLCELL_X1 FILLER_59_654 ();
 FILLCELL_X8 FILLER_59_690 ();
 FILLCELL_X4 FILLER_59_698 ();
 FILLCELL_X4 FILLER_59_722 ();
 FILLCELL_X2 FILLER_59_726 ();
 FILLCELL_X2 FILLER_59_742 ();
 FILLCELL_X1 FILLER_59_744 ();
 FILLCELL_X1 FILLER_59_750 ();
 FILLCELL_X2 FILLER_59_763 ();
 FILLCELL_X1 FILLER_59_765 ();
 FILLCELL_X4 FILLER_59_784 ();
 FILLCELL_X2 FILLER_59_788 ();
 FILLCELL_X4 FILLER_59_803 ();
 FILLCELL_X1 FILLER_59_807 ();
 FILLCELL_X2 FILLER_59_815 ();
 FILLCELL_X8 FILLER_59_833 ();
 FILLCELL_X4 FILLER_59_851 ();
 FILLCELL_X2 FILLER_59_855 ();
 FILLCELL_X8 FILLER_59_867 ();
 FILLCELL_X2 FILLER_59_875 ();
 FILLCELL_X1 FILLER_59_897 ();
 FILLCELL_X2 FILLER_59_922 ();
 FILLCELL_X8 FILLER_59_933 ();
 FILLCELL_X4 FILLER_59_941 ();
 FILLCELL_X2 FILLER_59_945 ();
 FILLCELL_X2 FILLER_59_975 ();
 FILLCELL_X2 FILLER_59_999 ();
 FILLCELL_X2 FILLER_59_1008 ();
 FILLCELL_X1 FILLER_59_1010 ();
 FILLCELL_X2 FILLER_59_1082 ();
 FILLCELL_X4 FILLER_59_1094 ();
 FILLCELL_X2 FILLER_59_1098 ();
 FILLCELL_X1 FILLER_59_1100 ();
 FILLCELL_X1 FILLER_59_1110 ();
 FILLCELL_X2 FILLER_59_1113 ();
 FILLCELL_X8 FILLER_59_1135 ();
 FILLCELL_X32 FILLER_59_1152 ();
 FILLCELL_X2 FILLER_59_1184 ();
 FILLCELL_X1 FILLER_59_1186 ();
 FILLCELL_X16 FILLER_59_1194 ();
 FILLCELL_X4 FILLER_59_1210 ();
 FILLCELL_X1 FILLER_59_1214 ();
 FILLCELL_X2 FILLER_59_1219 ();
 FILLCELL_X2 FILLER_59_1226 ();
 FILLCELL_X4 FILLER_60_17 ();
 FILLCELL_X2 FILLER_60_25 ();
 FILLCELL_X1 FILLER_60_27 ();
 FILLCELL_X32 FILLER_60_42 ();
 FILLCELL_X2 FILLER_60_74 ();
 FILLCELL_X1 FILLER_60_76 ();
 FILLCELL_X2 FILLER_60_84 ();
 FILLCELL_X16 FILLER_60_93 ();
 FILLCELL_X4 FILLER_60_109 ();
 FILLCELL_X1 FILLER_60_113 ();
 FILLCELL_X8 FILLER_60_116 ();
 FILLCELL_X2 FILLER_60_124 ();
 FILLCELL_X4 FILLER_60_133 ();
 FILLCELL_X1 FILLER_60_157 ();
 FILLCELL_X4 FILLER_60_165 ();
 FILLCELL_X2 FILLER_60_234 ();
 FILLCELL_X1 FILLER_60_249 ();
 FILLCELL_X1 FILLER_60_270 ();
 FILLCELL_X1 FILLER_60_278 ();
 FILLCELL_X2 FILLER_60_327 ();
 FILLCELL_X4 FILLER_60_334 ();
 FILLCELL_X4 FILLER_60_370 ();
 FILLCELL_X2 FILLER_60_374 ();
 FILLCELL_X4 FILLER_60_433 ();
 FILLCELL_X4 FILLER_60_457 ();
 FILLCELL_X1 FILLER_60_489 ();
 FILLCELL_X1 FILLER_60_503 ();
 FILLCELL_X1 FILLER_60_513 ();
 FILLCELL_X4 FILLER_60_524 ();
 FILLCELL_X1 FILLER_60_561 ();
 FILLCELL_X8 FILLER_60_571 ();
 FILLCELL_X2 FILLER_60_579 ();
 FILLCELL_X1 FILLER_60_581 ();
 FILLCELL_X4 FILLER_60_587 ();
 FILLCELL_X2 FILLER_60_591 ();
 FILLCELL_X1 FILLER_60_593 ();
 FILLCELL_X1 FILLER_60_607 ();
 FILLCELL_X4 FILLER_60_615 ();
 FILLCELL_X2 FILLER_60_619 ();
 FILLCELL_X2 FILLER_60_628 ();
 FILLCELL_X1 FILLER_60_630 ();
 FILLCELL_X4 FILLER_60_632 ();
 FILLCELL_X1 FILLER_60_636 ();
 FILLCELL_X4 FILLER_60_650 ();
 FILLCELL_X2 FILLER_60_678 ();
 FILLCELL_X8 FILLER_60_691 ();
 FILLCELL_X4 FILLER_60_699 ();
 FILLCELL_X2 FILLER_60_703 ();
 FILLCELL_X1 FILLER_60_705 ();
 FILLCELL_X4 FILLER_60_709 ();
 FILLCELL_X8 FILLER_60_729 ();
 FILLCELL_X16 FILLER_60_744 ();
 FILLCELL_X4 FILLER_60_760 ();
 FILLCELL_X8 FILLER_60_782 ();
 FILLCELL_X2 FILLER_60_790 ();
 FILLCELL_X1 FILLER_60_792 ();
 FILLCELL_X4 FILLER_60_807 ();
 FILLCELL_X1 FILLER_60_811 ();
 FILLCELL_X2 FILLER_60_819 ();
 FILLCELL_X1 FILLER_60_821 ();
 FILLCELL_X2 FILLER_60_833 ();
 FILLCELL_X1 FILLER_60_835 ();
 FILLCELL_X4 FILLER_60_853 ();
 FILLCELL_X1 FILLER_60_857 ();
 FILLCELL_X4 FILLER_60_872 ();
 FILLCELL_X4 FILLER_60_886 ();
 FILLCELL_X1 FILLER_60_890 ();
 FILLCELL_X8 FILLER_60_895 ();
 FILLCELL_X16 FILLER_60_934 ();
 FILLCELL_X8 FILLER_60_950 ();
 FILLCELL_X1 FILLER_60_958 ();
 FILLCELL_X4 FILLER_60_966 ();
 FILLCELL_X4 FILLER_60_974 ();
 FILLCELL_X8 FILLER_60_985 ();
 FILLCELL_X1 FILLER_60_993 ();
 FILLCELL_X8 FILLER_60_1021 ();
 FILLCELL_X4 FILLER_60_1029 ();
 FILLCELL_X2 FILLER_60_1033 ();
 FILLCELL_X8 FILLER_60_1044 ();
 FILLCELL_X1 FILLER_60_1052 ();
 FILLCELL_X4 FILLER_60_1056 ();
 FILLCELL_X4 FILLER_60_1062 ();
 FILLCELL_X8 FILLER_60_1069 ();
 FILLCELL_X2 FILLER_60_1077 ();
 FILLCELL_X1 FILLER_60_1079 ();
 FILLCELL_X16 FILLER_60_1085 ();
 FILLCELL_X2 FILLER_60_1101 ();
 FILLCELL_X1 FILLER_60_1189 ();
 FILLCELL_X2 FILLER_60_1201 ();
 FILLCELL_X2 FILLER_60_1210 ();
 FILLCELL_X1 FILLER_60_1212 ();
 FILLCELL_X8 FILLER_60_1240 ();
 FILLCELL_X4 FILLER_60_1248 ();
 FILLCELL_X2 FILLER_60_1252 ();
 FILLCELL_X1 FILLER_60_1254 ();
 FILLCELL_X2 FILLER_61_1 ();
 FILLCELL_X1 FILLER_61_3 ();
 FILLCELL_X4 FILLER_61_31 ();
 FILLCELL_X1 FILLER_61_35 ();
 FILLCELL_X8 FILLER_61_50 ();
 FILLCELL_X4 FILLER_61_58 ();
 FILLCELL_X1 FILLER_61_69 ();
 FILLCELL_X2 FILLER_61_77 ();
 FILLCELL_X2 FILLER_61_99 ();
 FILLCELL_X1 FILLER_61_101 ();
 FILLCELL_X1 FILLER_61_109 ();
 FILLCELL_X2 FILLER_61_130 ();
 FILLCELL_X1 FILLER_61_132 ();
 FILLCELL_X8 FILLER_61_167 ();
 FILLCELL_X4 FILLER_61_175 ();
 FILLCELL_X2 FILLER_61_179 ();
 FILLCELL_X1 FILLER_61_199 ();
 FILLCELL_X1 FILLER_61_223 ();
 FILLCELL_X1 FILLER_61_301 ();
 FILLCELL_X8 FILLER_61_316 ();
 FILLCELL_X4 FILLER_61_324 ();
 FILLCELL_X1 FILLER_61_328 ();
 FILLCELL_X8 FILLER_61_341 ();
 FILLCELL_X2 FILLER_61_354 ();
 FILLCELL_X8 FILLER_61_370 ();
 FILLCELL_X1 FILLER_61_378 ();
 FILLCELL_X2 FILLER_61_389 ();
 FILLCELL_X2 FILLER_61_411 ();
 FILLCELL_X4 FILLER_61_420 ();
 FILLCELL_X1 FILLER_61_445 ();
 FILLCELL_X2 FILLER_61_460 ();
 FILLCELL_X1 FILLER_61_462 ();
 FILLCELL_X4 FILLER_61_470 ();
 FILLCELL_X1 FILLER_61_474 ();
 FILLCELL_X8 FILLER_61_482 ();
 FILLCELL_X1 FILLER_61_490 ();
 FILLCELL_X8 FILLER_61_504 ();
 FILLCELL_X4 FILLER_61_519 ();
 FILLCELL_X2 FILLER_61_525 ();
 FILLCELL_X1 FILLER_61_527 ();
 FILLCELL_X2 FILLER_61_531 ();
 FILLCELL_X1 FILLER_61_533 ();
 FILLCELL_X8 FILLER_61_541 ();
 FILLCELL_X4 FILLER_61_549 ();
 FILLCELL_X1 FILLER_61_553 ();
 FILLCELL_X4 FILLER_61_558 ();
 FILLCELL_X2 FILLER_61_562 ();
 FILLCELL_X8 FILLER_61_588 ();
 FILLCELL_X2 FILLER_61_596 ();
 FILLCELL_X1 FILLER_61_598 ();
 FILLCELL_X2 FILLER_61_615 ();
 FILLCELL_X2 FILLER_61_631 ();
 FILLCELL_X1 FILLER_61_633 ();
 FILLCELL_X4 FILLER_61_641 ();
 FILLCELL_X4 FILLER_61_664 ();
 FILLCELL_X8 FILLER_61_673 ();
 FILLCELL_X2 FILLER_61_681 ();
 FILLCELL_X2 FILLER_61_696 ();
 FILLCELL_X2 FILLER_61_705 ();
 FILLCELL_X1 FILLER_61_707 ();
 FILLCELL_X16 FILLER_61_715 ();
 FILLCELL_X4 FILLER_61_731 ();
 FILLCELL_X1 FILLER_61_746 ();
 FILLCELL_X1 FILLER_61_751 ();
 FILLCELL_X1 FILLER_61_769 ();
 FILLCELL_X2 FILLER_61_772 ();
 FILLCELL_X2 FILLER_61_783 ();
 FILLCELL_X1 FILLER_61_785 ();
 FILLCELL_X2 FILLER_61_797 ();
 FILLCELL_X8 FILLER_61_802 ();
 FILLCELL_X4 FILLER_61_810 ();
 FILLCELL_X2 FILLER_61_814 ();
 FILLCELL_X1 FILLER_61_816 ();
 FILLCELL_X2 FILLER_61_827 ();
 FILLCELL_X4 FILLER_61_841 ();
 FILLCELL_X1 FILLER_61_845 ();
 FILLCELL_X2 FILLER_61_853 ();
 FILLCELL_X4 FILLER_61_872 ();
 FILLCELL_X2 FILLER_61_930 ();
 FILLCELL_X8 FILLER_61_939 ();
 FILLCELL_X2 FILLER_61_955 ();
 FILLCELL_X1 FILLER_61_957 ();
 FILLCELL_X2 FILLER_61_965 ();
 FILLCELL_X8 FILLER_61_981 ();
 FILLCELL_X4 FILLER_61_989 ();
 FILLCELL_X4 FILLER_61_997 ();
 FILLCELL_X2 FILLER_61_1001 ();
 FILLCELL_X4 FILLER_61_1009 ();
 FILLCELL_X2 FILLER_61_1051 ();
 FILLCELL_X4 FILLER_61_1060 ();
 FILLCELL_X2 FILLER_61_1064 ();
 FILLCELL_X8 FILLER_61_1095 ();
 FILLCELL_X4 FILLER_61_1103 ();
 FILLCELL_X2 FILLER_61_1107 ();
 FILLCELL_X4 FILLER_61_1132 ();
 FILLCELL_X4 FILLER_61_1150 ();
 FILLCELL_X1 FILLER_61_1154 ();
 FILLCELL_X8 FILLER_61_1172 ();
 FILLCELL_X2 FILLER_61_1180 ();
 FILLCELL_X2 FILLER_61_1220 ();
 FILLCELL_X1 FILLER_61_1222 ();
 FILLCELL_X8 FILLER_61_1245 ();
 FILLCELL_X2 FILLER_61_1253 ();
 FILLCELL_X2 FILLER_62_1 ();
 FILLCELL_X1 FILLER_62_3 ();
 FILLCELL_X2 FILLER_62_11 ();
 FILLCELL_X1 FILLER_62_13 ();
 FILLCELL_X4 FILLER_62_41 ();
 FILLCELL_X2 FILLER_62_45 ();
 FILLCELL_X1 FILLER_62_67 ();
 FILLCELL_X1 FILLER_62_88 ();
 FILLCELL_X1 FILLER_62_103 ();
 FILLCELL_X2 FILLER_62_138 ();
 FILLCELL_X1 FILLER_62_140 ();
 FILLCELL_X8 FILLER_62_155 ();
 FILLCELL_X4 FILLER_62_163 ();
 FILLCELL_X4 FILLER_62_204 ();
 FILLCELL_X2 FILLER_62_208 ();
 FILLCELL_X1 FILLER_62_243 ();
 FILLCELL_X2 FILLER_62_258 ();
 FILLCELL_X1 FILLER_62_260 ();
 FILLCELL_X1 FILLER_62_271 ();
 FILLCELL_X2 FILLER_62_318 ();
 FILLCELL_X1 FILLER_62_323 ();
 FILLCELL_X2 FILLER_62_337 ();
 FILLCELL_X4 FILLER_62_348 ();
 FILLCELL_X8 FILLER_62_355 ();
 FILLCELL_X4 FILLER_62_403 ();
 FILLCELL_X2 FILLER_62_407 ();
 FILLCELL_X1 FILLER_62_409 ();
 FILLCELL_X4 FILLER_62_435 ();
 FILLCELL_X1 FILLER_62_439 ();
 FILLCELL_X4 FILLER_62_447 ();
 FILLCELL_X16 FILLER_62_485 ();
 FILLCELL_X16 FILLER_62_514 ();
 FILLCELL_X4 FILLER_62_547 ();
 FILLCELL_X4 FILLER_62_560 ();
 FILLCELL_X2 FILLER_62_564 ();
 FILLCELL_X1 FILLER_62_566 ();
 FILLCELL_X4 FILLER_62_574 ();
 FILLCELL_X1 FILLER_62_578 ();
 FILLCELL_X4 FILLER_62_608 ();
 FILLCELL_X2 FILLER_62_612 ();
 FILLCELL_X1 FILLER_62_614 ();
 FILLCELL_X4 FILLER_62_626 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X2 FILLER_62_632 ();
 FILLCELL_X1 FILLER_62_634 ();
 FILLCELL_X8 FILLER_62_648 ();
 FILLCELL_X4 FILLER_62_656 ();
 FILLCELL_X2 FILLER_62_660 ();
 FILLCELL_X1 FILLER_62_662 ();
 FILLCELL_X2 FILLER_62_670 ();
 FILLCELL_X2 FILLER_62_675 ();
 FILLCELL_X1 FILLER_62_677 ();
 FILLCELL_X8 FILLER_62_691 ();
 FILLCELL_X2 FILLER_62_699 ();
 FILLCELL_X1 FILLER_62_701 ();
 FILLCELL_X1 FILLER_62_707 ();
 FILLCELL_X2 FILLER_62_724 ();
 FILLCELL_X2 FILLER_62_757 ();
 FILLCELL_X2 FILLER_62_777 ();
 FILLCELL_X1 FILLER_62_779 ();
 FILLCELL_X16 FILLER_62_793 ();
 FILLCELL_X8 FILLER_62_809 ();
 FILLCELL_X4 FILLER_62_829 ();
 FILLCELL_X1 FILLER_62_833 ();
 FILLCELL_X4 FILLER_62_836 ();
 FILLCELL_X8 FILLER_62_850 ();
 FILLCELL_X2 FILLER_62_858 ();
 FILLCELL_X4 FILLER_62_865 ();
 FILLCELL_X2 FILLER_62_869 ();
 FILLCELL_X16 FILLER_62_885 ();
 FILLCELL_X2 FILLER_62_901 ();
 FILLCELL_X4 FILLER_62_916 ();
 FILLCELL_X1 FILLER_62_969 ();
 FILLCELL_X1 FILLER_62_995 ();
 FILLCELL_X1 FILLER_62_1003 ();
 FILLCELL_X2 FILLER_62_1008 ();
 FILLCELL_X1 FILLER_62_1084 ();
 FILLCELL_X2 FILLER_62_1099 ();
 FILLCELL_X1 FILLER_62_1101 ();
 FILLCELL_X2 FILLER_62_1111 ();
 FILLCELL_X8 FILLER_62_1140 ();
 FILLCELL_X4 FILLER_62_1148 ();
 FILLCELL_X2 FILLER_62_1152 ();
 FILLCELL_X1 FILLER_62_1154 ();
 FILLCELL_X16 FILLER_62_1158 ();
 FILLCELL_X8 FILLER_62_1174 ();
 FILLCELL_X2 FILLER_62_1182 ();
 FILLCELL_X1 FILLER_62_1184 ();
 FILLCELL_X1 FILLER_62_1192 ();
 FILLCELL_X8 FILLER_62_1196 ();
 FILLCELL_X4 FILLER_62_1204 ();
 FILLCELL_X2 FILLER_62_1208 ();
 FILLCELL_X4 FILLER_62_1214 ();
 FILLCELL_X4 FILLER_62_1229 ();
 FILLCELL_X1 FILLER_62_1233 ();
 FILLCELL_X2 FILLER_62_1241 ();
 FILLCELL_X1 FILLER_62_1243 ();
 FILLCELL_X8 FILLER_62_1247 ();
 FILLCELL_X1 FILLER_63_1 ();
 FILLCELL_X2 FILLER_63_22 ();
 FILLCELL_X16 FILLER_63_45 ();
 FILLCELL_X1 FILLER_63_61 ();
 FILLCELL_X8 FILLER_63_70 ();
 FILLCELL_X2 FILLER_63_106 ();
 FILLCELL_X1 FILLER_63_108 ();
 FILLCELL_X4 FILLER_63_123 ();
 FILLCELL_X2 FILLER_63_127 ();
 FILLCELL_X1 FILLER_63_129 ();
 FILLCELL_X8 FILLER_63_144 ();
 FILLCELL_X4 FILLER_63_152 ();
 FILLCELL_X1 FILLER_63_193 ();
 FILLCELL_X4 FILLER_63_197 ();
 FILLCELL_X4 FILLER_63_208 ();
 FILLCELL_X2 FILLER_63_212 ();
 FILLCELL_X1 FILLER_63_214 ();
 FILLCELL_X2 FILLER_63_249 ();
 FILLCELL_X1 FILLER_63_251 ();
 FILLCELL_X1 FILLER_63_286 ();
 FILLCELL_X1 FILLER_63_290 ();
 FILLCELL_X2 FILLER_63_305 ();
 FILLCELL_X4 FILLER_63_327 ();
 FILLCELL_X2 FILLER_63_340 ();
 FILLCELL_X1 FILLER_63_342 ();
 FILLCELL_X4 FILLER_63_392 ();
 FILLCELL_X1 FILLER_63_396 ();
 FILLCELL_X16 FILLER_63_404 ();
 FILLCELL_X4 FILLER_63_420 ();
 FILLCELL_X2 FILLER_63_424 ();
 FILLCELL_X1 FILLER_63_426 ();
 FILLCELL_X4 FILLER_63_434 ();
 FILLCELL_X1 FILLER_63_438 ();
 FILLCELL_X16 FILLER_63_453 ();
 FILLCELL_X4 FILLER_63_469 ();
 FILLCELL_X1 FILLER_63_473 ();
 FILLCELL_X4 FILLER_63_501 ();
 FILLCELL_X2 FILLER_63_505 ();
 FILLCELL_X4 FILLER_63_537 ();
 FILLCELL_X8 FILLER_63_554 ();
 FILLCELL_X4 FILLER_63_569 ();
 FILLCELL_X2 FILLER_63_584 ();
 FILLCELL_X2 FILLER_63_604 ();
 FILLCELL_X1 FILLER_63_610 ();
 FILLCELL_X4 FILLER_63_630 ();
 FILLCELL_X2 FILLER_63_634 ();
 FILLCELL_X1 FILLER_63_636 ();
 FILLCELL_X2 FILLER_63_648 ();
 FILLCELL_X1 FILLER_63_650 ();
 FILLCELL_X2 FILLER_63_668 ();
 FILLCELL_X4 FILLER_63_674 ();
 FILLCELL_X4 FILLER_63_692 ();
 FILLCELL_X16 FILLER_63_701 ();
 FILLCELL_X8 FILLER_63_717 ();
 FILLCELL_X4 FILLER_63_743 ();
 FILLCELL_X1 FILLER_63_747 ();
 FILLCELL_X8 FILLER_63_753 ();
 FILLCELL_X1 FILLER_63_761 ();
 FILLCELL_X4 FILLER_63_774 ();
 FILLCELL_X2 FILLER_63_778 ();
 FILLCELL_X1 FILLER_63_787 ();
 FILLCELL_X2 FILLER_63_810 ();
 FILLCELL_X1 FILLER_63_812 ();
 FILLCELL_X8 FILLER_63_816 ();
 FILLCELL_X8 FILLER_63_827 ();
 FILLCELL_X4 FILLER_63_835 ();
 FILLCELL_X1 FILLER_63_839 ();
 FILLCELL_X4 FILLER_63_847 ();
 FILLCELL_X1 FILLER_63_851 ();
 FILLCELL_X2 FILLER_63_890 ();
 FILLCELL_X4 FILLER_63_904 ();
 FILLCELL_X2 FILLER_63_908 ();
 FILLCELL_X1 FILLER_63_910 ();
 FILLCELL_X8 FILLER_63_929 ();
 FILLCELL_X4 FILLER_63_943 ();
 FILLCELL_X16 FILLER_63_949 ();
 FILLCELL_X1 FILLER_63_965 ();
 FILLCELL_X1 FILLER_63_970 ();
 FILLCELL_X4 FILLER_63_974 ();
 FILLCELL_X2 FILLER_63_978 ();
 FILLCELL_X1 FILLER_63_980 ();
 FILLCELL_X4 FILLER_63_988 ();
 FILLCELL_X2 FILLER_63_992 ();
 FILLCELL_X2 FILLER_63_1009 ();
 FILLCELL_X1 FILLER_63_1011 ();
 FILLCELL_X4 FILLER_63_1016 ();
 FILLCELL_X2 FILLER_63_1027 ();
 FILLCELL_X1 FILLER_63_1037 ();
 FILLCELL_X2 FILLER_63_1041 ();
 FILLCELL_X4 FILLER_63_1070 ();
 FILLCELL_X2 FILLER_63_1074 ();
 FILLCELL_X1 FILLER_63_1076 ();
 FILLCELL_X8 FILLER_63_1104 ();
 FILLCELL_X2 FILLER_63_1112 ();
 FILLCELL_X2 FILLER_63_1162 ();
 FILLCELL_X1 FILLER_63_1164 ();
 FILLCELL_X4 FILLER_63_1187 ();
 FILLCELL_X1 FILLER_63_1191 ();
 FILLCELL_X2 FILLER_63_1212 ();
 FILLCELL_X4 FILLER_63_1218 ();
 FILLCELL_X1 FILLER_63_1222 ();
 FILLCELL_X4 FILLER_63_1228 ();
 FILLCELL_X2 FILLER_63_1232 ();
 FILLCELL_X1 FILLER_63_1234 ();
 FILLCELL_X16 FILLER_64_1 ();
 FILLCELL_X4 FILLER_64_17 ();
 FILLCELL_X4 FILLER_64_42 ();
 FILLCELL_X2 FILLER_64_46 ();
 FILLCELL_X1 FILLER_64_48 ();
 FILLCELL_X4 FILLER_64_76 ();
 FILLCELL_X1 FILLER_64_80 ();
 FILLCELL_X2 FILLER_64_88 ();
 FILLCELL_X1 FILLER_64_90 ();
 FILLCELL_X4 FILLER_64_98 ();
 FILLCELL_X4 FILLER_64_129 ();
 FILLCELL_X1 FILLER_64_133 ();
 FILLCELL_X4 FILLER_64_139 ();
 FILLCELL_X1 FILLER_64_143 ();
 FILLCELL_X4 FILLER_64_192 ();
 FILLCELL_X1 FILLER_64_196 ();
 FILLCELL_X2 FILLER_64_211 ();
 FILLCELL_X1 FILLER_64_213 ();
 FILLCELL_X4 FILLER_64_221 ();
 FILLCELL_X4 FILLER_64_248 ();
 FILLCELL_X1 FILLER_64_252 ();
 FILLCELL_X4 FILLER_64_273 ();
 FILLCELL_X1 FILLER_64_277 ();
 FILLCELL_X2 FILLER_64_291 ();
 FILLCELL_X1 FILLER_64_293 ();
 FILLCELL_X1 FILLER_64_298 ();
 FILLCELL_X1 FILLER_64_302 ();
 FILLCELL_X2 FILLER_64_310 ();
 FILLCELL_X1 FILLER_64_312 ();
 FILLCELL_X4 FILLER_64_316 ();
 FILLCELL_X1 FILLER_64_322 ();
 FILLCELL_X2 FILLER_64_350 ();
 FILLCELL_X2 FILLER_64_377 ();
 FILLCELL_X1 FILLER_64_379 ();
 FILLCELL_X1 FILLER_64_401 ();
 FILLCELL_X4 FILLER_64_412 ();
 FILLCELL_X8 FILLER_64_423 ();
 FILLCELL_X1 FILLER_64_431 ();
 FILLCELL_X8 FILLER_64_436 ();
 FILLCELL_X4 FILLER_64_447 ();
 FILLCELL_X4 FILLER_64_458 ();
 FILLCELL_X4 FILLER_64_465 ();
 FILLCELL_X2 FILLER_64_469 ();
 FILLCELL_X1 FILLER_64_471 ();
 FILLCELL_X1 FILLER_64_476 ();
 FILLCELL_X8 FILLER_64_480 ();
 FILLCELL_X2 FILLER_64_488 ();
 FILLCELL_X4 FILLER_64_517 ();
 FILLCELL_X2 FILLER_64_521 ();
 FILLCELL_X1 FILLER_64_523 ();
 FILLCELL_X1 FILLER_64_537 ();
 FILLCELL_X8 FILLER_64_545 ();
 FILLCELL_X4 FILLER_64_553 ();
 FILLCELL_X1 FILLER_64_557 ();
 FILLCELL_X2 FILLER_64_577 ();
 FILLCELL_X8 FILLER_64_586 ();
 FILLCELL_X2 FILLER_64_594 ();
 FILLCELL_X2 FILLER_64_620 ();
 FILLCELL_X1 FILLER_64_643 ();
 FILLCELL_X2 FILLER_64_653 ();
 FILLCELL_X1 FILLER_64_655 ();
 FILLCELL_X4 FILLER_64_674 ();
 FILLCELL_X2 FILLER_64_685 ();
 FILLCELL_X8 FILLER_64_698 ();
 FILLCELL_X4 FILLER_64_706 ();
 FILLCELL_X2 FILLER_64_710 ();
 FILLCELL_X1 FILLER_64_712 ();
 FILLCELL_X16 FILLER_64_723 ();
 FILLCELL_X4 FILLER_64_739 ();
 FILLCELL_X2 FILLER_64_743 ();
 FILLCELL_X1 FILLER_64_745 ();
 FILLCELL_X16 FILLER_64_776 ();
 FILLCELL_X2 FILLER_64_792 ();
 FILLCELL_X8 FILLER_64_797 ();
 FILLCELL_X4 FILLER_64_805 ();
 FILLCELL_X2 FILLER_64_809 ();
 FILLCELL_X2 FILLER_64_837 ();
 FILLCELL_X4 FILLER_64_856 ();
 FILLCELL_X2 FILLER_64_865 ();
 FILLCELL_X1 FILLER_64_867 ();
 FILLCELL_X2 FILLER_64_875 ();
 FILLCELL_X2 FILLER_64_881 ();
 FILLCELL_X2 FILLER_64_892 ();
 FILLCELL_X1 FILLER_64_935 ();
 FILLCELL_X4 FILLER_64_956 ();
 FILLCELL_X2 FILLER_64_960 ();
 FILLCELL_X8 FILLER_64_976 ();
 FILLCELL_X4 FILLER_64_984 ();
 FILLCELL_X2 FILLER_64_988 ();
 FILLCELL_X8 FILLER_64_997 ();
 FILLCELL_X1 FILLER_64_1005 ();
 FILLCELL_X1 FILLER_64_1044 ();
 FILLCELL_X1 FILLER_64_1049 ();
 FILLCELL_X1 FILLER_64_1060 ();
 FILLCELL_X16 FILLER_64_1083 ();
 FILLCELL_X2 FILLER_64_1099 ();
 FILLCELL_X1 FILLER_64_1106 ();
 FILLCELL_X4 FILLER_64_1112 ();
 FILLCELL_X1 FILLER_64_1116 ();
 FILLCELL_X8 FILLER_64_1136 ();
 FILLCELL_X4 FILLER_64_1144 ();
 FILLCELL_X1 FILLER_64_1148 ();
 FILLCELL_X1 FILLER_64_1155 ();
 FILLCELL_X1 FILLER_64_1167 ();
 FILLCELL_X1 FILLER_64_1182 ();
 FILLCELL_X1 FILLER_64_1192 ();
 FILLCELL_X1 FILLER_64_1196 ();
 FILLCELL_X1 FILLER_64_1204 ();
 FILLCELL_X1 FILLER_64_1212 ();
 FILLCELL_X1 FILLER_64_1218 ();
 FILLCELL_X4 FILLER_64_1224 ();
 FILLCELL_X2 FILLER_65_1 ();
 FILLCELL_X2 FILLER_65_10 ();
 FILLCELL_X8 FILLER_65_39 ();
 FILLCELL_X4 FILLER_65_47 ();
 FILLCELL_X1 FILLER_65_51 ();
 FILLCELL_X4 FILLER_65_59 ();
 FILLCELL_X1 FILLER_65_63 ();
 FILLCELL_X4 FILLER_65_91 ();
 FILLCELL_X2 FILLER_65_115 ();
 FILLCELL_X1 FILLER_65_117 ();
 FILLCELL_X4 FILLER_65_132 ();
 FILLCELL_X1 FILLER_65_136 ();
 FILLCELL_X8 FILLER_65_176 ();
 FILLCELL_X4 FILLER_65_198 ();
 FILLCELL_X2 FILLER_65_202 ();
 FILLCELL_X2 FILLER_65_215 ();
 FILLCELL_X1 FILLER_65_217 ();
 FILLCELL_X1 FILLER_65_239 ();
 FILLCELL_X4 FILLER_65_251 ();
 FILLCELL_X2 FILLER_65_255 ();
 FILLCELL_X1 FILLER_65_257 ();
 FILLCELL_X1 FILLER_65_262 ();
 FILLCELL_X8 FILLER_65_266 ();
 FILLCELL_X2 FILLER_65_333 ();
 FILLCELL_X1 FILLER_65_335 ();
 FILLCELL_X4 FILLER_65_363 ();
 FILLCELL_X2 FILLER_65_374 ();
 FILLCELL_X1 FILLER_65_376 ();
 FILLCELL_X2 FILLER_65_487 ();
 FILLCELL_X1 FILLER_65_489 ();
 FILLCELL_X1 FILLER_65_535 ();
 FILLCELL_X16 FILLER_65_553 ();
 FILLCELL_X1 FILLER_65_569 ();
 FILLCELL_X8 FILLER_65_584 ();
 FILLCELL_X2 FILLER_65_592 ();
 FILLCELL_X2 FILLER_65_607 ();
 FILLCELL_X1 FILLER_65_609 ();
 FILLCELL_X2 FILLER_65_619 ();
 FILLCELL_X4 FILLER_65_625 ();
 FILLCELL_X4 FILLER_65_640 ();
 FILLCELL_X2 FILLER_65_647 ();
 FILLCELL_X2 FILLER_65_690 ();
 FILLCELL_X1 FILLER_65_692 ();
 FILLCELL_X1 FILLER_65_716 ();
 FILLCELL_X1 FILLER_65_724 ();
 FILLCELL_X2 FILLER_65_738 ();
 FILLCELL_X2 FILLER_65_759 ();
 FILLCELL_X2 FILLER_65_772 ();
 FILLCELL_X2 FILLER_65_791 ();
 FILLCELL_X8 FILLER_65_813 ();
 FILLCELL_X4 FILLER_65_821 ();
 FILLCELL_X8 FILLER_65_828 ();
 FILLCELL_X4 FILLER_65_843 ();
 FILLCELL_X2 FILLER_65_847 ();
 FILLCELL_X1 FILLER_65_849 ();
 FILLCELL_X4 FILLER_65_867 ();
 FILLCELL_X1 FILLER_65_871 ();
 FILLCELL_X8 FILLER_65_906 ();
 FILLCELL_X2 FILLER_65_914 ();
 FILLCELL_X2 FILLER_65_923 ();
 FILLCELL_X16 FILLER_65_929 ();
 FILLCELL_X4 FILLER_65_947 ();
 FILLCELL_X4 FILLER_65_976 ();
 FILLCELL_X2 FILLER_65_980 ();
 FILLCELL_X4 FILLER_65_989 ();
 FILLCELL_X2 FILLER_65_993 ();
 FILLCELL_X1 FILLER_65_995 ();
 FILLCELL_X2 FILLER_65_1006 ();
 FILLCELL_X1 FILLER_65_1008 ();
 FILLCELL_X8 FILLER_65_1021 ();
 FILLCELL_X8 FILLER_65_1033 ();
 FILLCELL_X1 FILLER_65_1041 ();
 FILLCELL_X8 FILLER_65_1073 ();
 FILLCELL_X4 FILLER_65_1081 ();
 FILLCELL_X1 FILLER_65_1085 ();
 FILLCELL_X8 FILLER_65_1108 ();
 FILLCELL_X2 FILLER_65_1147 ();
 FILLCELL_X4 FILLER_65_1171 ();
 FILLCELL_X2 FILLER_65_1175 ();
 FILLCELL_X1 FILLER_65_1177 ();
 FILLCELL_X4 FILLER_65_1198 ();
 FILLCELL_X1 FILLER_65_1202 ();
 FILLCELL_X8 FILLER_65_1243 ();
 FILLCELL_X4 FILLER_65_1251 ();
 FILLCELL_X2 FILLER_66_26 ();
 FILLCELL_X1 FILLER_66_28 ();
 FILLCELL_X4 FILLER_66_50 ();
 FILLCELL_X2 FILLER_66_54 ();
 FILLCELL_X2 FILLER_66_97 ();
 FILLCELL_X1 FILLER_66_106 ();
 FILLCELL_X4 FILLER_66_114 ();
 FILLCELL_X4 FILLER_66_139 ();
 FILLCELL_X1 FILLER_66_143 ();
 FILLCELL_X16 FILLER_66_153 ();
 FILLCELL_X8 FILLER_66_169 ();
 FILLCELL_X4 FILLER_66_177 ();
 FILLCELL_X4 FILLER_66_201 ();
 FILLCELL_X2 FILLER_66_205 ();
 FILLCELL_X1 FILLER_66_214 ();
 FILLCELL_X4 FILLER_66_293 ();
 FILLCELL_X2 FILLER_66_297 ();
 FILLCELL_X2 FILLER_66_322 ();
 FILLCELL_X2 FILLER_66_345 ();
 FILLCELL_X1 FILLER_66_347 ();
 FILLCELL_X4 FILLER_66_355 ();
 FILLCELL_X2 FILLER_66_359 ();
 FILLCELL_X1 FILLER_66_361 ();
 FILLCELL_X1 FILLER_66_389 ();
 FILLCELL_X1 FILLER_66_428 ();
 FILLCELL_X2 FILLER_66_450 ();
 FILLCELL_X1 FILLER_66_452 ();
 FILLCELL_X1 FILLER_66_461 ();
 FILLCELL_X32 FILLER_66_493 ();
 FILLCELL_X8 FILLER_66_525 ();
 FILLCELL_X1 FILLER_66_533 ();
 FILLCELL_X2 FILLER_66_547 ();
 FILLCELL_X8 FILLER_66_562 ();
 FILLCELL_X4 FILLER_66_594 ();
 FILLCELL_X2 FILLER_66_603 ();
 FILLCELL_X2 FILLER_66_622 ();
 FILLCELL_X4 FILLER_66_650 ();
 FILLCELL_X4 FILLER_66_667 ();
 FILLCELL_X1 FILLER_66_678 ();
 FILLCELL_X2 FILLER_66_706 ();
 FILLCELL_X1 FILLER_66_708 ();
 FILLCELL_X4 FILLER_66_723 ();
 FILLCELL_X2 FILLER_66_727 ();
 FILLCELL_X2 FILLER_66_736 ();
 FILLCELL_X4 FILLER_66_747 ();
 FILLCELL_X1 FILLER_66_751 ();
 FILLCELL_X8 FILLER_66_763 ();
 FILLCELL_X2 FILLER_66_771 ();
 FILLCELL_X4 FILLER_66_784 ();
 FILLCELL_X1 FILLER_66_788 ();
 FILLCELL_X4 FILLER_66_797 ();
 FILLCELL_X2 FILLER_66_801 ();
 FILLCELL_X1 FILLER_66_803 ();
 FILLCELL_X16 FILLER_66_828 ();
 FILLCELL_X2 FILLER_66_844 ();
 FILLCELL_X8 FILLER_66_853 ();
 FILLCELL_X8 FILLER_66_870 ();
 FILLCELL_X2 FILLER_66_878 ();
 FILLCELL_X4 FILLER_66_883 ();
 FILLCELL_X1 FILLER_66_887 ();
 FILLCELL_X4 FILLER_66_892 ();
 FILLCELL_X2 FILLER_66_896 ();
 FILLCELL_X1 FILLER_66_898 ();
 FILLCELL_X1 FILLER_66_906 ();
 FILLCELL_X8 FILLER_66_940 ();
 FILLCELL_X2 FILLER_66_948 ();
 FILLCELL_X4 FILLER_66_952 ();
 FILLCELL_X2 FILLER_66_956 ();
 FILLCELL_X8 FILLER_66_972 ();
 FILLCELL_X4 FILLER_66_987 ();
 FILLCELL_X1 FILLER_66_991 ();
 FILLCELL_X4 FILLER_66_1014 ();
 FILLCELL_X4 FILLER_66_1047 ();
 FILLCELL_X2 FILLER_66_1051 ();
 FILLCELL_X1 FILLER_66_1053 ();
 FILLCELL_X2 FILLER_66_1061 ();
 FILLCELL_X16 FILLER_66_1096 ();
 FILLCELL_X1 FILLER_66_1112 ();
 FILLCELL_X8 FILLER_66_1125 ();
 FILLCELL_X4 FILLER_66_1133 ();
 FILLCELL_X2 FILLER_66_1137 ();
 FILLCELL_X1 FILLER_66_1139 ();
 FILLCELL_X4 FILLER_66_1142 ();
 FILLCELL_X2 FILLER_66_1146 ();
 FILLCELL_X1 FILLER_66_1148 ();
 FILLCELL_X2 FILLER_66_1152 ();
 FILLCELL_X1 FILLER_66_1154 ();
 FILLCELL_X4 FILLER_66_1207 ();
 FILLCELL_X2 FILLER_66_1211 ();
 FILLCELL_X4 FILLER_66_1217 ();
 FILLCELL_X1 FILLER_66_1221 ();
 FILLCELL_X16 FILLER_66_1226 ();
 FILLCELL_X2 FILLER_66_1242 ();
 FILLCELL_X1 FILLER_66_1244 ();
 FILLCELL_X2 FILLER_66_1253 ();
 FILLCELL_X4 FILLER_67_1 ();
 FILLCELL_X1 FILLER_67_5 ();
 FILLCELL_X4 FILLER_67_33 ();
 FILLCELL_X1 FILLER_67_37 ();
 FILLCELL_X2 FILLER_67_45 ();
 FILLCELL_X2 FILLER_67_54 ();
 FILLCELL_X1 FILLER_67_56 ();
 FILLCELL_X8 FILLER_67_84 ();
 FILLCELL_X4 FILLER_67_92 ();
 FILLCELL_X2 FILLER_67_96 ();
 FILLCELL_X4 FILLER_67_125 ();
 FILLCELL_X1 FILLER_67_129 ();
 FILLCELL_X8 FILLER_67_137 ();
 FILLCELL_X1 FILLER_67_145 ();
 FILLCELL_X4 FILLER_67_153 ();
 FILLCELL_X1 FILLER_67_157 ();
 FILLCELL_X4 FILLER_67_205 ();
 FILLCELL_X2 FILLER_67_213 ();
 FILLCELL_X1 FILLER_67_215 ();
 FILLCELL_X4 FILLER_67_223 ();
 FILLCELL_X8 FILLER_67_248 ();
 FILLCELL_X4 FILLER_67_256 ();
 FILLCELL_X8 FILLER_67_276 ();
 FILLCELL_X4 FILLER_67_284 ();
 FILLCELL_X1 FILLER_67_288 ();
 FILLCELL_X1 FILLER_67_316 ();
 FILLCELL_X2 FILLER_67_330 ();
 FILLCELL_X4 FILLER_67_347 ();
 FILLCELL_X4 FILLER_67_360 ();
 FILLCELL_X1 FILLER_67_408 ();
 FILLCELL_X2 FILLER_67_419 ();
 FILLCELL_X1 FILLER_67_421 ();
 FILLCELL_X4 FILLER_67_425 ();
 FILLCELL_X1 FILLER_67_436 ();
 FILLCELL_X1 FILLER_67_444 ();
 FILLCELL_X2 FILLER_67_472 ();
 FILLCELL_X1 FILLER_67_474 ();
 FILLCELL_X1 FILLER_67_478 ();
 FILLCELL_X2 FILLER_67_499 ();
 FILLCELL_X1 FILLER_67_501 ();
 FILLCELL_X16 FILLER_67_509 ();
 FILLCELL_X2 FILLER_67_525 ();
 FILLCELL_X1 FILLER_67_527 ();
 FILLCELL_X16 FILLER_67_545 ();
 FILLCELL_X2 FILLER_67_561 ();
 FILLCELL_X2 FILLER_67_580 ();
 FILLCELL_X1 FILLER_67_582 ();
 FILLCELL_X1 FILLER_67_585 ();
 FILLCELL_X8 FILLER_67_593 ();
 FILLCELL_X2 FILLER_67_601 ();
 FILLCELL_X2 FILLER_67_630 ();
 FILLCELL_X1 FILLER_67_632 ();
 FILLCELL_X16 FILLER_67_635 ();
 FILLCELL_X8 FILLER_67_651 ();
 FILLCELL_X1 FILLER_67_659 ();
 FILLCELL_X16 FILLER_67_689 ();
 FILLCELL_X8 FILLER_67_705 ();
 FILLCELL_X2 FILLER_67_713 ();
 FILLCELL_X8 FILLER_67_722 ();
 FILLCELL_X2 FILLER_67_730 ();
 FILLCELL_X8 FILLER_67_766 ();
 FILLCELL_X4 FILLER_67_816 ();
 FILLCELL_X1 FILLER_67_823 ();
 FILLCELL_X4 FILLER_67_831 ();
 FILLCELL_X4 FILLER_67_842 ();
 FILLCELL_X2 FILLER_67_846 ();
 FILLCELL_X1 FILLER_67_848 ();
 FILLCELL_X2 FILLER_67_851 ();
 FILLCELL_X1 FILLER_67_853 ();
 FILLCELL_X8 FILLER_67_871 ();
 FILLCELL_X2 FILLER_67_879 ();
 FILLCELL_X1 FILLER_67_881 ();
 FILLCELL_X16 FILLER_67_892 ();
 FILLCELL_X8 FILLER_67_908 ();
 FILLCELL_X1 FILLER_67_916 ();
 FILLCELL_X4 FILLER_67_924 ();
 FILLCELL_X1 FILLER_67_928 ();
 FILLCELL_X8 FILLER_67_946 ();
 FILLCELL_X2 FILLER_67_954 ();
 FILLCELL_X1 FILLER_67_956 ();
 FILLCELL_X2 FILLER_67_968 ();
 FILLCELL_X4 FILLER_67_976 ();
 FILLCELL_X8 FILLER_67_1029 ();
 FILLCELL_X2 FILLER_67_1037 ();
 FILLCELL_X1 FILLER_67_1039 ();
 FILLCELL_X16 FILLER_67_1045 ();
 FILLCELL_X8 FILLER_67_1061 ();
 FILLCELL_X2 FILLER_67_1086 ();
 FILLCELL_X1 FILLER_67_1088 ();
 FILLCELL_X2 FILLER_67_1093 ();
 FILLCELL_X4 FILLER_67_1097 ();
 FILLCELL_X1 FILLER_67_1101 ();
 FILLCELL_X2 FILLER_67_1105 ();
 FILLCELL_X4 FILLER_67_1129 ();
 FILLCELL_X2 FILLER_67_1133 ();
 FILLCELL_X4 FILLER_67_1161 ();
 FILLCELL_X1 FILLER_67_1165 ();
 FILLCELL_X1 FILLER_67_1168 ();
 FILLCELL_X2 FILLER_67_1198 ();
 FILLCELL_X4 FILLER_67_1203 ();
 FILLCELL_X1 FILLER_67_1207 ();
 FILLCELL_X4 FILLER_67_1217 ();
 FILLCELL_X2 FILLER_67_1221 ();
 FILLCELL_X8 FILLER_68_1 ();
 FILLCELL_X2 FILLER_68_9 ();
 FILLCELL_X1 FILLER_68_11 ();
 FILLCELL_X2 FILLER_68_39 ();
 FILLCELL_X1 FILLER_68_41 ();
 FILLCELL_X16 FILLER_68_49 ();
 FILLCELL_X8 FILLER_68_65 ();
 FILLCELL_X4 FILLER_68_73 ();
 FILLCELL_X2 FILLER_68_77 ();
 FILLCELL_X8 FILLER_68_98 ();
 FILLCELL_X2 FILLER_68_127 ();
 FILLCELL_X1 FILLER_68_129 ();
 FILLCELL_X16 FILLER_68_164 ();
 FILLCELL_X4 FILLER_68_180 ();
 FILLCELL_X2 FILLER_68_184 ();
 FILLCELL_X4 FILLER_68_251 ();
 FILLCELL_X2 FILLER_68_255 ();
 FILLCELL_X2 FILLER_68_282 ();
 FILLCELL_X1 FILLER_68_284 ();
 FILLCELL_X2 FILLER_68_292 ();
 FILLCELL_X1 FILLER_68_294 ();
 FILLCELL_X2 FILLER_68_308 ();
 FILLCELL_X1 FILLER_68_310 ();
 FILLCELL_X2 FILLER_68_398 ();
 FILLCELL_X1 FILLER_68_400 ();
 FILLCELL_X2 FILLER_68_414 ();
 FILLCELL_X8 FILLER_68_446 ();
 FILLCELL_X2 FILLER_68_454 ();
 FILLCELL_X2 FILLER_68_466 ();
 FILLCELL_X4 FILLER_68_479 ();
 FILLCELL_X2 FILLER_68_483 ();
 FILLCELL_X1 FILLER_68_489 ();
 FILLCELL_X1 FILLER_68_493 ();
 FILLCELL_X16 FILLER_68_521 ();
 FILLCELL_X16 FILLER_68_556 ();
 FILLCELL_X8 FILLER_68_572 ();
 FILLCELL_X4 FILLER_68_580 ();
 FILLCELL_X1 FILLER_68_591 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X4 FILLER_68_632 ();
 FILLCELL_X8 FILLER_68_670 ();
 FILLCELL_X2 FILLER_68_678 ();
 FILLCELL_X2 FILLER_68_688 ();
 FILLCELL_X4 FILLER_68_710 ();
 FILLCELL_X2 FILLER_68_714 ();
 FILLCELL_X8 FILLER_68_723 ();
 FILLCELL_X4 FILLER_68_731 ();
 FILLCELL_X1 FILLER_68_735 ();
 FILLCELL_X2 FILLER_68_745 ();
 FILLCELL_X2 FILLER_68_765 ();
 FILLCELL_X1 FILLER_68_767 ();
 FILLCELL_X8 FILLER_68_772 ();
 FILLCELL_X1 FILLER_68_794 ();
 FILLCELL_X8 FILLER_68_802 ();
 FILLCELL_X1 FILLER_68_817 ();
 FILLCELL_X1 FILLER_68_825 ();
 FILLCELL_X4 FILLER_68_833 ();
 FILLCELL_X2 FILLER_68_837 ();
 FILLCELL_X1 FILLER_68_839 ();
 FILLCELL_X16 FILLER_68_847 ();
 FILLCELL_X8 FILLER_68_863 ();
 FILLCELL_X4 FILLER_68_871 ();
 FILLCELL_X2 FILLER_68_875 ();
 FILLCELL_X1 FILLER_68_937 ();
 FILLCELL_X2 FILLER_68_941 ();
 FILLCELL_X2 FILLER_68_956 ();
 FILLCELL_X4 FILLER_68_978 ();
 FILLCELL_X2 FILLER_68_982 ();
 FILLCELL_X1 FILLER_68_984 ();
 FILLCELL_X8 FILLER_68_996 ();
 FILLCELL_X4 FILLER_68_1004 ();
 FILLCELL_X2 FILLER_68_1008 ();
 FILLCELL_X1 FILLER_68_1041 ();
 FILLCELL_X8 FILLER_68_1046 ();
 FILLCELL_X2 FILLER_68_1054 ();
 FILLCELL_X1 FILLER_68_1056 ();
 FILLCELL_X4 FILLER_68_1064 ();
 FILLCELL_X2 FILLER_68_1078 ();
 FILLCELL_X1 FILLER_68_1080 ();
 FILLCELL_X2 FILLER_68_1119 ();
 FILLCELL_X1 FILLER_68_1121 ();
 FILLCELL_X2 FILLER_68_1130 ();
 FILLCELL_X4 FILLER_68_1138 ();
 FILLCELL_X16 FILLER_68_1176 ();
 FILLCELL_X4 FILLER_68_1192 ();
 FILLCELL_X1 FILLER_68_1232 ();
 FILLCELL_X16 FILLER_68_1236 ();
 FILLCELL_X2 FILLER_68_1252 ();
 FILLCELL_X1 FILLER_68_1254 ();
 FILLCELL_X16 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_17 ();
 FILLCELL_X1 FILLER_69_21 ();
 FILLCELL_X4 FILLER_69_29 ();
 FILLCELL_X1 FILLER_69_33 ();
 FILLCELL_X4 FILLER_69_41 ();
 FILLCELL_X2 FILLER_69_45 ();
 FILLCELL_X8 FILLER_69_54 ();
 FILLCELL_X2 FILLER_69_62 ();
 FILLCELL_X4 FILLER_69_71 ();
 FILLCELL_X2 FILLER_69_75 ();
 FILLCELL_X4 FILLER_69_84 ();
 FILLCELL_X4 FILLER_69_129 ();
 FILLCELL_X1 FILLER_69_140 ();
 FILLCELL_X8 FILLER_69_150 ();
 FILLCELL_X2 FILLER_69_158 ();
 FILLCELL_X1 FILLER_69_160 ();
 FILLCELL_X16 FILLER_69_193 ();
 FILLCELL_X8 FILLER_69_209 ();
 FILLCELL_X4 FILLER_69_217 ();
 FILLCELL_X2 FILLER_69_221 ();
 FILLCELL_X1 FILLER_69_223 ();
 FILLCELL_X4 FILLER_69_330 ();
 FILLCELL_X2 FILLER_69_334 ();
 FILLCELL_X1 FILLER_69_341 ();
 FILLCELL_X1 FILLER_69_351 ();
 FILLCELL_X1 FILLER_69_362 ();
 FILLCELL_X4 FILLER_69_370 ();
 FILLCELL_X2 FILLER_69_374 ();
 FILLCELL_X1 FILLER_69_376 ();
 FILLCELL_X2 FILLER_69_384 ();
 FILLCELL_X1 FILLER_69_390 ();
 FILLCELL_X8 FILLER_69_401 ();
 FILLCELL_X4 FILLER_69_409 ();
 FILLCELL_X1 FILLER_69_433 ();
 FILLCELL_X1 FILLER_69_441 ();
 FILLCELL_X1 FILLER_69_462 ();
 FILLCELL_X1 FILLER_69_477 ();
 FILLCELL_X8 FILLER_69_485 ();
 FILLCELL_X1 FILLER_69_493 ();
 FILLCELL_X8 FILLER_69_501 ();
 FILLCELL_X1 FILLER_69_509 ();
 FILLCELL_X4 FILLER_69_537 ();
 FILLCELL_X2 FILLER_69_541 ();
 FILLCELL_X2 FILLER_69_546 ();
 FILLCELL_X1 FILLER_69_548 ();
 FILLCELL_X2 FILLER_69_562 ();
 FILLCELL_X1 FILLER_69_564 ();
 FILLCELL_X4 FILLER_69_591 ();
 FILLCELL_X2 FILLER_69_595 ();
 FILLCELL_X1 FILLER_69_597 ();
 FILLCELL_X2 FILLER_69_605 ();
 FILLCELL_X1 FILLER_69_607 ();
 FILLCELL_X1 FILLER_69_621 ();
 FILLCELL_X2 FILLER_69_624 ();
 FILLCELL_X4 FILLER_69_635 ();
 FILLCELL_X1 FILLER_69_639 ();
 FILLCELL_X2 FILLER_69_643 ();
 FILLCELL_X1 FILLER_69_650 ();
 FILLCELL_X8 FILLER_69_681 ();
 FILLCELL_X2 FILLER_69_689 ();
 FILLCELL_X2 FILLER_69_705 ();
 FILLCELL_X1 FILLER_69_707 ();
 FILLCELL_X2 FILLER_69_715 ();
 FILLCELL_X1 FILLER_69_717 ();
 FILLCELL_X2 FILLER_69_725 ();
 FILLCELL_X1 FILLER_69_727 ();
 FILLCELL_X2 FILLER_69_737 ();
 FILLCELL_X1 FILLER_69_739 ();
 FILLCELL_X2 FILLER_69_756 ();
 FILLCELL_X1 FILLER_69_809 ();
 FILLCELL_X16 FILLER_69_817 ();
 FILLCELL_X4 FILLER_69_833 ();
 FILLCELL_X1 FILLER_69_837 ();
 FILLCELL_X4 FILLER_69_841 ();
 FILLCELL_X2 FILLER_69_845 ();
 FILLCELL_X1 FILLER_69_847 ();
 FILLCELL_X4 FILLER_69_855 ();
 FILLCELL_X1 FILLER_69_859 ();
 FILLCELL_X1 FILLER_69_874 ();
 FILLCELL_X1 FILLER_69_878 ();
 FILLCELL_X1 FILLER_69_896 ();
 FILLCELL_X16 FILLER_69_913 ();
 FILLCELL_X1 FILLER_69_946 ();
 FILLCELL_X4 FILLER_69_954 ();
 FILLCELL_X16 FILLER_69_967 ();
 FILLCELL_X8 FILLER_69_983 ();
 FILLCELL_X1 FILLER_69_998 ();
 FILLCELL_X8 FILLER_69_1023 ();
 FILLCELL_X4 FILLER_69_1031 ();
 FILLCELL_X1 FILLER_69_1035 ();
 FILLCELL_X8 FILLER_69_1044 ();
 FILLCELL_X1 FILLER_69_1052 ();
 FILLCELL_X2 FILLER_69_1073 ();
 FILLCELL_X2 FILLER_69_1097 ();
 FILLCELL_X1 FILLER_69_1131 ();
 FILLCELL_X4 FILLER_69_1154 ();
 FILLCELL_X1 FILLER_69_1158 ();
 FILLCELL_X4 FILLER_69_1166 ();
 FILLCELL_X1 FILLER_69_1170 ();
 FILLCELL_X4 FILLER_69_1178 ();
 FILLCELL_X1 FILLER_69_1192 ();
 FILLCELL_X8 FILLER_69_1207 ();
 FILLCELL_X2 FILLER_69_1215 ();
 FILLCELL_X4 FILLER_69_1224 ();
 FILLCELL_X2 FILLER_69_1228 ();
 FILLCELL_X1 FILLER_69_1230 ();
 FILLCELL_X2 FILLER_69_1253 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X4 FILLER_70_12 ();
 FILLCELL_X2 FILLER_70_16 ();
 FILLCELL_X1 FILLER_70_18 ();
 FILLCELL_X1 FILLER_70_46 ();
 FILLCELL_X1 FILLER_70_108 ();
 FILLCELL_X4 FILLER_70_116 ();
 FILLCELL_X8 FILLER_70_127 ();
 FILLCELL_X4 FILLER_70_135 ();
 FILLCELL_X2 FILLER_70_139 ();
 FILLCELL_X1 FILLER_70_141 ();
 FILLCELL_X1 FILLER_70_149 ();
 FILLCELL_X8 FILLER_70_183 ();
 FILLCELL_X4 FILLER_70_191 ();
 FILLCELL_X1 FILLER_70_195 ();
 FILLCELL_X4 FILLER_70_208 ();
 FILLCELL_X1 FILLER_70_212 ();
 FILLCELL_X2 FILLER_70_253 ();
 FILLCELL_X16 FILLER_70_328 ();
 FILLCELL_X4 FILLER_70_344 ();
 FILLCELL_X1 FILLER_70_348 ();
 FILLCELL_X1 FILLER_70_354 ();
 FILLCELL_X1 FILLER_70_367 ();
 FILLCELL_X1 FILLER_70_379 ();
 FILLCELL_X1 FILLER_70_404 ();
 FILLCELL_X8 FILLER_70_412 ();
 FILLCELL_X4 FILLER_70_420 ();
 FILLCELL_X1 FILLER_70_473 ();
 FILLCELL_X2 FILLER_70_494 ();
 FILLCELL_X2 FILLER_70_499 ();
 FILLCELL_X2 FILLER_70_505 ();
 FILLCELL_X8 FILLER_70_517 ();
 FILLCELL_X1 FILLER_70_525 ();
 FILLCELL_X2 FILLER_70_539 ();
 FILLCELL_X1 FILLER_70_541 ();
 FILLCELL_X2 FILLER_70_558 ();
 FILLCELL_X8 FILLER_70_567 ();
 FILLCELL_X4 FILLER_70_575 ();
 FILLCELL_X1 FILLER_70_579 ();
 FILLCELL_X8 FILLER_70_587 ();
 FILLCELL_X2 FILLER_70_595 ();
 FILLCELL_X4 FILLER_70_604 ();
 FILLCELL_X1 FILLER_70_608 ();
 FILLCELL_X16 FILLER_70_612 ();
 FILLCELL_X2 FILLER_70_628 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X1 FILLER_70_632 ();
 FILLCELL_X1 FILLER_70_636 ();
 FILLCELL_X2 FILLER_70_649 ();
 FILLCELL_X1 FILLER_70_651 ();
 FILLCELL_X1 FILLER_70_654 ();
 FILLCELL_X2 FILLER_70_659 ();
 FILLCELL_X1 FILLER_70_661 ();
 FILLCELL_X2 FILLER_70_665 ();
 FILLCELL_X2 FILLER_70_672 ();
 FILLCELL_X8 FILLER_70_681 ();
 FILLCELL_X4 FILLER_70_689 ();
 FILLCELL_X2 FILLER_70_693 ();
 FILLCELL_X1 FILLER_70_695 ();
 FILLCELL_X2 FILLER_70_713 ();
 FILLCELL_X1 FILLER_70_715 ();
 FILLCELL_X1 FILLER_70_719 ();
 FILLCELL_X1 FILLER_70_724 ();
 FILLCELL_X1 FILLER_70_728 ();
 FILLCELL_X1 FILLER_70_743 ();
 FILLCELL_X2 FILLER_70_758 ();
 FILLCELL_X1 FILLER_70_760 ();
 FILLCELL_X2 FILLER_70_770 ();
 FILLCELL_X1 FILLER_70_772 ();
 FILLCELL_X2 FILLER_70_802 ();
 FILLCELL_X1 FILLER_70_804 ();
 FILLCELL_X2 FILLER_70_826 ();
 FILLCELL_X2 FILLER_70_835 ();
 FILLCELL_X1 FILLER_70_837 ();
 FILLCELL_X4 FILLER_70_845 ();
 FILLCELL_X1 FILLER_70_849 ();
 FILLCELL_X1 FILLER_70_864 ();
 FILLCELL_X8 FILLER_70_868 ();
 FILLCELL_X4 FILLER_70_883 ();
 FILLCELL_X1 FILLER_70_887 ();
 FILLCELL_X1 FILLER_70_891 ();
 FILLCELL_X2 FILLER_70_899 ();
 FILLCELL_X1 FILLER_70_939 ();
 FILLCELL_X4 FILLER_70_943 ();
 FILLCELL_X1 FILLER_70_947 ();
 FILLCELL_X4 FILLER_70_970 ();
 FILLCELL_X1 FILLER_70_974 ();
 FILLCELL_X4 FILLER_70_982 ();
 FILLCELL_X8 FILLER_70_988 ();
 FILLCELL_X4 FILLER_70_996 ();
 FILLCELL_X1 FILLER_70_1000 ();
 FILLCELL_X2 FILLER_70_1003 ();
 FILLCELL_X1 FILLER_70_1012 ();
 FILLCELL_X2 FILLER_70_1045 ();
 FILLCELL_X4 FILLER_70_1062 ();
 FILLCELL_X2 FILLER_70_1066 ();
 FILLCELL_X1 FILLER_70_1075 ();
 FILLCELL_X8 FILLER_70_1079 ();
 FILLCELL_X2 FILLER_70_1087 ();
 FILLCELL_X1 FILLER_70_1089 ();
 FILLCELL_X1 FILLER_70_1094 ();
 FILLCELL_X4 FILLER_70_1120 ();
 FILLCELL_X1 FILLER_70_1138 ();
 FILLCELL_X8 FILLER_70_1145 ();
 FILLCELL_X1 FILLER_70_1153 ();
 FILLCELL_X8 FILLER_70_1157 ();
 FILLCELL_X1 FILLER_70_1165 ();
 FILLCELL_X8 FILLER_70_1177 ();
 FILLCELL_X16 FILLER_70_1192 ();
 FILLCELL_X1 FILLER_70_1208 ();
 FILLCELL_X4 FILLER_70_1216 ();
 FILLCELL_X1 FILLER_70_1220 ();
 FILLCELL_X8 FILLER_70_1224 ();
 FILLCELL_X1 FILLER_70_1232 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X4 FILLER_71_25 ();
 FILLCELL_X2 FILLER_71_29 ();
 FILLCELL_X1 FILLER_71_31 ();
 FILLCELL_X4 FILLER_71_39 ();
 FILLCELL_X1 FILLER_71_43 ();
 FILLCELL_X1 FILLER_71_58 ();
 FILLCELL_X1 FILLER_71_66 ();
 FILLCELL_X2 FILLER_71_87 ();
 FILLCELL_X1 FILLER_71_89 ();
 FILLCELL_X4 FILLER_71_104 ();
 FILLCELL_X2 FILLER_71_128 ();
 FILLCELL_X4 FILLER_71_150 ();
 FILLCELL_X8 FILLER_71_190 ();
 FILLCELL_X8 FILLER_71_205 ();
 FILLCELL_X2 FILLER_71_213 ();
 FILLCELL_X1 FILLER_71_215 ();
 FILLCELL_X4 FILLER_71_223 ();
 FILLCELL_X1 FILLER_71_231 ();
 FILLCELL_X4 FILLER_71_258 ();
 FILLCELL_X1 FILLER_71_262 ();
 FILLCELL_X2 FILLER_71_284 ();
 FILLCELL_X1 FILLER_71_286 ();
 FILLCELL_X1 FILLER_71_307 ();
 FILLCELL_X1 FILLER_71_328 ();
 FILLCELL_X4 FILLER_71_334 ();
 FILLCELL_X8 FILLER_71_345 ();
 FILLCELL_X2 FILLER_71_353 ();
 FILLCELL_X1 FILLER_71_355 ();
 FILLCELL_X4 FILLER_71_392 ();
 FILLCELL_X1 FILLER_71_396 ();
 FILLCELL_X1 FILLER_71_404 ();
 FILLCELL_X1 FILLER_71_436 ();
 FILLCELL_X2 FILLER_71_440 ();
 FILLCELL_X1 FILLER_71_449 ();
 FILLCELL_X2 FILLER_71_454 ();
 FILLCELL_X1 FILLER_71_477 ();
 FILLCELL_X2 FILLER_71_498 ();
 FILLCELL_X2 FILLER_71_520 ();
 FILLCELL_X1 FILLER_71_522 ();
 FILLCELL_X16 FILLER_71_530 ();
 FILLCELL_X4 FILLER_71_553 ();
 FILLCELL_X2 FILLER_71_557 ();
 FILLCELL_X1 FILLER_71_595 ();
 FILLCELL_X2 FILLER_71_613 ();
 FILLCELL_X2 FILLER_71_619 ();
 FILLCELL_X2 FILLER_71_626 ();
 FILLCELL_X2 FILLER_71_637 ();
 FILLCELL_X4 FILLER_71_659 ();
 FILLCELL_X1 FILLER_71_663 ();
 FILLCELL_X16 FILLER_71_676 ();
 FILLCELL_X8 FILLER_71_692 ();
 FILLCELL_X4 FILLER_71_700 ();
 FILLCELL_X2 FILLER_71_704 ();
 FILLCELL_X1 FILLER_71_706 ();
 FILLCELL_X1 FILLER_71_714 ();
 FILLCELL_X1 FILLER_71_720 ();
 FILLCELL_X1 FILLER_71_725 ();
 FILLCELL_X2 FILLER_71_730 ();
 FILLCELL_X2 FILLER_71_740 ();
 FILLCELL_X1 FILLER_71_742 ();
 FILLCELL_X2 FILLER_71_748 ();
 FILLCELL_X1 FILLER_71_750 ();
 FILLCELL_X2 FILLER_71_756 ();
 FILLCELL_X1 FILLER_71_758 ();
 FILLCELL_X4 FILLER_71_784 ();
 FILLCELL_X2 FILLER_71_788 ();
 FILLCELL_X1 FILLER_71_790 ();
 FILLCELL_X2 FILLER_71_812 ();
 FILLCELL_X1 FILLER_71_814 ();
 FILLCELL_X2 FILLER_71_831 ();
 FILLCELL_X1 FILLER_71_833 ();
 FILLCELL_X8 FILLER_71_841 ();
 FILLCELL_X1 FILLER_71_849 ();
 FILLCELL_X8 FILLER_71_867 ();
 FILLCELL_X2 FILLER_71_882 ();
 FILLCELL_X2 FILLER_71_891 ();
 FILLCELL_X16 FILLER_71_916 ();
 FILLCELL_X2 FILLER_71_932 ();
 FILLCELL_X1 FILLER_71_934 ();
 FILLCELL_X1 FILLER_71_947 ();
 FILLCELL_X2 FILLER_71_955 ();
 FILLCELL_X1 FILLER_71_957 ();
 FILLCELL_X1 FILLER_71_960 ();
 FILLCELL_X16 FILLER_71_988 ();
 FILLCELL_X1 FILLER_71_1004 ();
 FILLCELL_X2 FILLER_71_1008 ();
 FILLCELL_X1 FILLER_71_1010 ();
 FILLCELL_X4 FILLER_71_1021 ();
 FILLCELL_X2 FILLER_71_1025 ();
 FILLCELL_X1 FILLER_71_1027 ();
 FILLCELL_X8 FILLER_71_1035 ();
 FILLCELL_X4 FILLER_71_1066 ();
 FILLCELL_X1 FILLER_71_1070 ();
 FILLCELL_X8 FILLER_71_1104 ();
 FILLCELL_X4 FILLER_71_1112 ();
 FILLCELL_X2 FILLER_71_1116 ();
 FILLCELL_X1 FILLER_71_1118 ();
 FILLCELL_X2 FILLER_71_1123 ();
 FILLCELL_X1 FILLER_71_1125 ();
 FILLCELL_X2 FILLER_71_1132 ();
 FILLCELL_X1 FILLER_71_1134 ();
 FILLCELL_X4 FILLER_71_1162 ();
 FILLCELL_X8 FILLER_71_1180 ();
 FILLCELL_X2 FILLER_71_1210 ();
 FILLCELL_X4 FILLER_71_1232 ();
 FILLCELL_X1 FILLER_71_1236 ();
 FILLCELL_X4 FILLER_71_1244 ();
 FILLCELL_X2 FILLER_71_1248 ();
 FILLCELL_X1 FILLER_71_1250 ();
 FILLCELL_X8 FILLER_72_1 ();
 FILLCELL_X2 FILLER_72_9 ();
 FILLCELL_X2 FILLER_72_38 ();
 FILLCELL_X1 FILLER_72_40 ();
 FILLCELL_X4 FILLER_72_61 ();
 FILLCELL_X2 FILLER_72_85 ();
 FILLCELL_X1 FILLER_72_87 ();
 FILLCELL_X8 FILLER_72_102 ();
 FILLCELL_X4 FILLER_72_110 ();
 FILLCELL_X2 FILLER_72_114 ();
 FILLCELL_X1 FILLER_72_116 ();
 FILLCELL_X4 FILLER_72_151 ();
 FILLCELL_X1 FILLER_72_155 ();
 FILLCELL_X4 FILLER_72_163 ();
 FILLCELL_X1 FILLER_72_167 ();
 FILLCELL_X2 FILLER_72_187 ();
 FILLCELL_X1 FILLER_72_189 ();
 FILLCELL_X1 FILLER_72_210 ();
 FILLCELL_X1 FILLER_72_221 ();
 FILLCELL_X1 FILLER_72_265 ();
 FILLCELL_X8 FILLER_72_273 ();
 FILLCELL_X4 FILLER_72_281 ();
 FILLCELL_X1 FILLER_72_293 ();
 FILLCELL_X1 FILLER_72_307 ();
 FILLCELL_X8 FILLER_72_345 ();
 FILLCELL_X1 FILLER_72_353 ();
 FILLCELL_X2 FILLER_72_379 ();
 FILLCELL_X1 FILLER_72_381 ();
 FILLCELL_X2 FILLER_72_420 ();
 FILLCELL_X1 FILLER_72_429 ();
 FILLCELL_X4 FILLER_72_450 ();
 FILLCELL_X1 FILLER_72_454 ();
 FILLCELL_X1 FILLER_72_469 ();
 FILLCELL_X4 FILLER_72_477 ();
 FILLCELL_X2 FILLER_72_481 ();
 FILLCELL_X2 FILLER_72_510 ();
 FILLCELL_X4 FILLER_72_519 ();
 FILLCELL_X2 FILLER_72_523 ();
 FILLCELL_X1 FILLER_72_525 ();
 FILLCELL_X8 FILLER_72_535 ();
 FILLCELL_X2 FILLER_72_543 ();
 FILLCELL_X32 FILLER_72_558 ();
 FILLCELL_X2 FILLER_72_590 ();
 FILLCELL_X2 FILLER_72_599 ();
 FILLCELL_X2 FILLER_72_608 ();
 FILLCELL_X1 FILLER_72_610 ();
 FILLCELL_X4 FILLER_72_615 ();
 FILLCELL_X1 FILLER_72_641 ();
 FILLCELL_X2 FILLER_72_666 ();
 FILLCELL_X16 FILLER_72_683 ();
 FILLCELL_X4 FILLER_72_699 ();
 FILLCELL_X2 FILLER_72_703 ();
 FILLCELL_X1 FILLER_72_708 ();
 FILLCELL_X2 FILLER_72_721 ();
 FILLCELL_X2 FILLER_72_727 ();
 FILLCELL_X1 FILLER_72_729 ();
 FILLCELL_X2 FILLER_72_737 ();
 FILLCELL_X1 FILLER_72_739 ();
 FILLCELL_X1 FILLER_72_744 ();
 FILLCELL_X4 FILLER_72_749 ();
 FILLCELL_X2 FILLER_72_753 ();
 FILLCELL_X1 FILLER_72_755 ();
 FILLCELL_X1 FILLER_72_778 ();
 FILLCELL_X1 FILLER_72_782 ();
 FILLCELL_X2 FILLER_72_790 ();
 FILLCELL_X2 FILLER_72_825 ();
 FILLCELL_X1 FILLER_72_827 ();
 FILLCELL_X1 FILLER_72_835 ();
 FILLCELL_X1 FILLER_72_843 ();
 FILLCELL_X1 FILLER_72_851 ();
 FILLCELL_X2 FILLER_72_859 ();
 FILLCELL_X4 FILLER_72_875 ();
 FILLCELL_X8 FILLER_72_896 ();
 FILLCELL_X4 FILLER_72_904 ();
 FILLCELL_X1 FILLER_72_908 ();
 FILLCELL_X1 FILLER_72_929 ();
 FILLCELL_X8 FILLER_72_972 ();
 FILLCELL_X2 FILLER_72_980 ();
 FILLCELL_X4 FILLER_72_999 ();
 FILLCELL_X1 FILLER_72_1003 ();
 FILLCELL_X8 FILLER_72_1010 ();
 FILLCELL_X8 FILLER_72_1021 ();
 FILLCELL_X1 FILLER_72_1029 ();
 FILLCELL_X8 FILLER_72_1050 ();
 FILLCELL_X1 FILLER_72_1058 ();
 FILLCELL_X4 FILLER_72_1115 ();
 FILLCELL_X2 FILLER_72_1129 ();
 FILLCELL_X8 FILLER_72_1153 ();
 FILLCELL_X1 FILLER_72_1161 ();
 FILLCELL_X2 FILLER_72_1168 ();
 FILLCELL_X1 FILLER_72_1170 ();
 FILLCELL_X4 FILLER_72_1218 ();
 FILLCELL_X2 FILLER_72_1222 ();
 FILLCELL_X1 FILLER_72_1234 ();
 FILLCELL_X1 FILLER_73_1 ();
 FILLCELL_X1 FILLER_73_9 ();
 FILLCELL_X1 FILLER_73_37 ();
 FILLCELL_X16 FILLER_73_45 ();
 FILLCELL_X2 FILLER_73_61 ();
 FILLCELL_X8 FILLER_73_97 ();
 FILLCELL_X2 FILLER_73_105 ();
 FILLCELL_X1 FILLER_73_107 ();
 FILLCELL_X2 FILLER_73_115 ();
 FILLCELL_X1 FILLER_73_117 ();
 FILLCELL_X4 FILLER_73_125 ();
 FILLCELL_X2 FILLER_73_129 ();
 FILLCELL_X1 FILLER_73_131 ();
 FILLCELL_X2 FILLER_73_139 ();
 FILLCELL_X1 FILLER_73_155 ();
 FILLCELL_X4 FILLER_73_164 ();
 FILLCELL_X2 FILLER_73_168 ();
 FILLCELL_X1 FILLER_73_170 ();
 FILLCELL_X4 FILLER_73_177 ();
 FILLCELL_X1 FILLER_73_192 ();
 FILLCELL_X8 FILLER_73_200 ();
 FILLCELL_X4 FILLER_73_208 ();
 FILLCELL_X2 FILLER_73_236 ();
 FILLCELL_X1 FILLER_73_265 ();
 FILLCELL_X4 FILLER_73_276 ();
 FILLCELL_X2 FILLER_73_280 ();
 FILLCELL_X4 FILLER_73_308 ();
 FILLCELL_X4 FILLER_73_362 ();
 FILLCELL_X2 FILLER_73_366 ();
 FILLCELL_X2 FILLER_73_375 ();
 FILLCELL_X1 FILLER_73_377 ();
 FILLCELL_X2 FILLER_73_382 ();
 FILLCELL_X1 FILLER_73_384 ();
 FILLCELL_X16 FILLER_73_388 ();
 FILLCELL_X8 FILLER_73_404 ();
 FILLCELL_X8 FILLER_73_415 ();
 FILLCELL_X4 FILLER_73_427 ();
 FILLCELL_X4 FILLER_73_451 ();
 FILLCELL_X1 FILLER_73_455 ();
 FILLCELL_X4 FILLER_73_464 ();
 FILLCELL_X1 FILLER_73_473 ();
 FILLCELL_X4 FILLER_73_477 ();
 FILLCELL_X2 FILLER_73_481 ();
 FILLCELL_X2 FILLER_73_490 ();
 FILLCELL_X1 FILLER_73_492 ();
 FILLCELL_X16 FILLER_73_507 ();
 FILLCELL_X8 FILLER_73_523 ();
 FILLCELL_X1 FILLER_73_531 ();
 FILLCELL_X1 FILLER_73_536 ();
 FILLCELL_X16 FILLER_73_540 ();
 FILLCELL_X8 FILLER_73_556 ();
 FILLCELL_X1 FILLER_73_564 ();
 FILLCELL_X2 FILLER_73_583 ();
 FILLCELL_X1 FILLER_73_585 ();
 FILLCELL_X8 FILLER_73_604 ();
 FILLCELL_X1 FILLER_73_612 ();
 FILLCELL_X8 FILLER_73_681 ();
 FILLCELL_X2 FILLER_73_689 ();
 FILLCELL_X1 FILLER_73_691 ();
 FILLCELL_X2 FILLER_73_699 ();
 FILLCELL_X1 FILLER_73_701 ();
 FILLCELL_X2 FILLER_73_711 ();
 FILLCELL_X1 FILLER_73_713 ();
 FILLCELL_X2 FILLER_73_721 ();
 FILLCELL_X1 FILLER_73_727 ();
 FILLCELL_X2 FILLER_73_733 ();
 FILLCELL_X4 FILLER_73_753 ();
 FILLCELL_X4 FILLER_73_762 ();
 FILLCELL_X2 FILLER_73_766 ();
 FILLCELL_X1 FILLER_73_768 ();
 FILLCELL_X2 FILLER_73_773 ();
 FILLCELL_X4 FILLER_73_788 ();
 FILLCELL_X4 FILLER_73_796 ();
 FILLCELL_X2 FILLER_73_812 ();
 FILLCELL_X1 FILLER_73_814 ();
 FILLCELL_X1 FILLER_73_822 ();
 FILLCELL_X1 FILLER_73_837 ();
 FILLCELL_X4 FILLER_73_849 ();
 FILLCELL_X32 FILLER_73_858 ();
 FILLCELL_X4 FILLER_73_931 ();
 FILLCELL_X8 FILLER_73_950 ();
 FILLCELL_X2 FILLER_73_958 ();
 FILLCELL_X1 FILLER_73_960 ();
 FILLCELL_X4 FILLER_73_968 ();
 FILLCELL_X8 FILLER_73_987 ();
 FILLCELL_X2 FILLER_73_995 ();
 FILLCELL_X16 FILLER_73_1018 ();
 FILLCELL_X4 FILLER_73_1034 ();
 FILLCELL_X2 FILLER_73_1038 ();
 FILLCELL_X1 FILLER_73_1047 ();
 FILLCELL_X8 FILLER_73_1052 ();
 FILLCELL_X2 FILLER_73_1060 ();
 FILLCELL_X1 FILLER_73_1062 ();
 FILLCELL_X8 FILLER_73_1068 ();
 FILLCELL_X2 FILLER_73_1076 ();
 FILLCELL_X1 FILLER_73_1078 ();
 FILLCELL_X8 FILLER_73_1090 ();
 FILLCELL_X4 FILLER_73_1098 ();
 FILLCELL_X1 FILLER_73_1102 ();
 FILLCELL_X8 FILLER_73_1124 ();
 FILLCELL_X4 FILLER_73_1132 ();
 FILLCELL_X2 FILLER_73_1136 ();
 FILLCELL_X1 FILLER_73_1138 ();
 FILLCELL_X4 FILLER_73_1150 ();
 FILLCELL_X1 FILLER_73_1154 ();
 FILLCELL_X8 FILLER_73_1172 ();
 FILLCELL_X4 FILLER_73_1180 ();
 FILLCELL_X2 FILLER_73_1184 ();
 FILLCELL_X1 FILLER_73_1189 ();
 FILLCELL_X1 FILLER_73_1202 ();
 FILLCELL_X4 FILLER_73_1223 ();
 FILLCELL_X2 FILLER_73_1227 ();
 FILLCELL_X1 FILLER_73_1229 ();
 FILLCELL_X4 FILLER_73_1250 ();
 FILLCELL_X1 FILLER_73_1254 ();
 FILLCELL_X4 FILLER_74_1 ();
 FILLCELL_X16 FILLER_74_46 ();
 FILLCELL_X4 FILLER_74_62 ();
 FILLCELL_X2 FILLER_74_66 ();
 FILLCELL_X1 FILLER_74_68 ();
 FILLCELL_X4 FILLER_74_76 ();
 FILLCELL_X4 FILLER_74_94 ();
 FILLCELL_X1 FILLER_74_98 ();
 FILLCELL_X16 FILLER_74_106 ();
 FILLCELL_X4 FILLER_74_122 ();
 FILLCELL_X1 FILLER_74_126 ();
 FILLCELL_X2 FILLER_74_134 ();
 FILLCELL_X1 FILLER_74_143 ();
 FILLCELL_X1 FILLER_74_147 ();
 FILLCELL_X1 FILLER_74_155 ();
 FILLCELL_X8 FILLER_74_166 ();
 FILLCELL_X1 FILLER_74_177 ();
 FILLCELL_X2 FILLER_74_185 ();
 FILLCELL_X2 FILLER_74_207 ();
 FILLCELL_X1 FILLER_74_209 ();
 FILLCELL_X1 FILLER_74_217 ();
 FILLCELL_X1 FILLER_74_230 ();
 FILLCELL_X2 FILLER_74_241 ();
 FILLCELL_X1 FILLER_74_243 ();
 FILLCELL_X4 FILLER_74_251 ();
 FILLCELL_X1 FILLER_74_255 ();
 FILLCELL_X2 FILLER_74_263 ();
 FILLCELL_X2 FILLER_74_272 ();
 FILLCELL_X1 FILLER_74_274 ();
 FILLCELL_X2 FILLER_74_278 ();
 FILLCELL_X1 FILLER_74_280 ();
 FILLCELL_X4 FILLER_74_288 ();
 FILLCELL_X2 FILLER_74_292 ();
 FILLCELL_X2 FILLER_74_298 ();
 FILLCELL_X8 FILLER_74_303 ();
 FILLCELL_X2 FILLER_74_315 ();
 FILLCELL_X1 FILLER_74_317 ();
 FILLCELL_X2 FILLER_74_321 ();
 FILLCELL_X4 FILLER_74_330 ();
 FILLCELL_X2 FILLER_74_334 ();
 FILLCELL_X1 FILLER_74_336 ();
 FILLCELL_X4 FILLER_74_357 ();
 FILLCELL_X1 FILLER_74_361 ();
 FILLCELL_X8 FILLER_74_403 ();
 FILLCELL_X4 FILLER_74_411 ();
 FILLCELL_X4 FILLER_74_419 ();
 FILLCELL_X16 FILLER_74_426 ();
 FILLCELL_X4 FILLER_74_442 ();
 FILLCELL_X2 FILLER_74_458 ();
 FILLCELL_X1 FILLER_74_472 ();
 FILLCELL_X2 FILLER_74_489 ();
 FILLCELL_X2 FILLER_74_563 ();
 FILLCELL_X1 FILLER_74_565 ();
 FILLCELL_X16 FILLER_74_573 ();
 FILLCELL_X2 FILLER_74_589 ();
 FILLCELL_X1 FILLER_74_591 ();
 FILLCELL_X2 FILLER_74_658 ();
 FILLCELL_X16 FILLER_74_684 ();
 FILLCELL_X4 FILLER_74_700 ();
 FILLCELL_X2 FILLER_74_704 ();
 FILLCELL_X2 FILLER_74_716 ();
 FILLCELL_X2 FILLER_74_722 ();
 FILLCELL_X1 FILLER_74_724 ();
 FILLCELL_X16 FILLER_74_729 ();
 FILLCELL_X4 FILLER_74_745 ();
 FILLCELL_X1 FILLER_74_749 ();
 FILLCELL_X16 FILLER_74_757 ();
 FILLCELL_X1 FILLER_74_773 ();
 FILLCELL_X4 FILLER_74_788 ();
 FILLCELL_X4 FILLER_74_831 ();
 FILLCELL_X2 FILLER_74_835 ();
 FILLCELL_X1 FILLER_74_837 ();
 FILLCELL_X1 FILLER_74_842 ();
 FILLCELL_X2 FILLER_74_850 ();
 FILLCELL_X4 FILLER_74_866 ();
 FILLCELL_X16 FILLER_74_877 ();
 FILLCELL_X4 FILLER_74_893 ();
 FILLCELL_X2 FILLER_74_897 ();
 FILLCELL_X4 FILLER_74_926 ();
 FILLCELL_X2 FILLER_74_930 ();
 FILLCELL_X1 FILLER_74_932 ();
 FILLCELL_X2 FILLER_74_958 ();
 FILLCELL_X1 FILLER_74_960 ();
 FILLCELL_X8 FILLER_74_983 ();
 FILLCELL_X2 FILLER_74_991 ();
 FILLCELL_X1 FILLER_74_993 ();
 FILLCELL_X4 FILLER_74_1000 ();
 FILLCELL_X2 FILLER_74_1004 ();
 FILLCELL_X1 FILLER_74_1063 ();
 FILLCELL_X8 FILLER_74_1068 ();
 FILLCELL_X1 FILLER_74_1076 ();
 FILLCELL_X1 FILLER_74_1087 ();
 FILLCELL_X4 FILLER_74_1099 ();
 FILLCELL_X4 FILLER_74_1114 ();
 FILLCELL_X1 FILLER_74_1118 ();
 FILLCELL_X2 FILLER_74_1121 ();
 FILLCELL_X8 FILLER_74_1133 ();
 FILLCELL_X4 FILLER_74_1141 ();
 FILLCELL_X1 FILLER_74_1145 ();
 FILLCELL_X2 FILLER_74_1160 ();
 FILLCELL_X1 FILLER_74_1162 ();
 FILLCELL_X8 FILLER_74_1167 ();
 FILLCELL_X2 FILLER_74_1175 ();
 FILLCELL_X1 FILLER_74_1202 ();
 FILLCELL_X1 FILLER_74_1231 ();
 FILLCELL_X2 FILLER_74_1235 ();
 FILLCELL_X1 FILLER_74_1237 ();
 FILLCELL_X8 FILLER_74_1244 ();
 FILLCELL_X16 FILLER_75_1 ();
 FILLCELL_X4 FILLER_75_17 ();
 FILLCELL_X8 FILLER_75_36 ();
 FILLCELL_X4 FILLER_75_44 ();
 FILLCELL_X1 FILLER_75_95 ();
 FILLCELL_X1 FILLER_75_103 ();
 FILLCELL_X8 FILLER_75_111 ();
 FILLCELL_X1 FILLER_75_119 ();
 FILLCELL_X4 FILLER_75_140 ();
 FILLCELL_X2 FILLER_75_144 ();
 FILLCELL_X8 FILLER_75_149 ();
 FILLCELL_X1 FILLER_75_157 ();
 FILLCELL_X2 FILLER_75_178 ();
 FILLCELL_X1 FILLER_75_180 ();
 FILLCELL_X2 FILLER_75_186 ();
 FILLCELL_X1 FILLER_75_188 ();
 FILLCELL_X4 FILLER_75_196 ();
 FILLCELL_X1 FILLER_75_207 ();
 FILLCELL_X2 FILLER_75_228 ();
 FILLCELL_X4 FILLER_75_244 ();
 FILLCELL_X2 FILLER_75_248 ();
 FILLCELL_X4 FILLER_75_257 ();
 FILLCELL_X2 FILLER_75_261 ();
 FILLCELL_X1 FILLER_75_263 ();
 FILLCELL_X4 FILLER_75_277 ();
 FILLCELL_X1 FILLER_75_281 ();
 FILLCELL_X2 FILLER_75_302 ();
 FILLCELL_X1 FILLER_75_304 ();
 FILLCELL_X4 FILLER_75_325 ();
 FILLCELL_X4 FILLER_75_369 ();
 FILLCELL_X1 FILLER_75_373 ();
 FILLCELL_X4 FILLER_75_384 ();
 FILLCELL_X1 FILLER_75_388 ();
 FILLCELL_X1 FILLER_75_399 ();
 FILLCELL_X1 FILLER_75_409 ();
 FILLCELL_X1 FILLER_75_419 ();
 FILLCELL_X4 FILLER_75_427 ();
 FILLCELL_X1 FILLER_75_435 ();
 FILLCELL_X2 FILLER_75_439 ();
 FILLCELL_X1 FILLER_75_441 ();
 FILLCELL_X1 FILLER_75_481 ();
 FILLCELL_X2 FILLER_75_489 ();
 FILLCELL_X1 FILLER_75_491 ();
 FILLCELL_X4 FILLER_75_521 ();
 FILLCELL_X1 FILLER_75_525 ();
 FILLCELL_X4 FILLER_75_552 ();
 FILLCELL_X2 FILLER_75_556 ();
 FILLCELL_X1 FILLER_75_558 ();
 FILLCELL_X32 FILLER_75_566 ();
 FILLCELL_X4 FILLER_75_598 ();
 FILLCELL_X1 FILLER_75_602 ();
 FILLCELL_X4 FILLER_75_608 ();
 FILLCELL_X2 FILLER_75_612 ();
 FILLCELL_X2 FILLER_75_621 ();
 FILLCELL_X2 FILLER_75_661 ();
 FILLCELL_X2 FILLER_75_679 ();
 FILLCELL_X4 FILLER_75_690 ();
 FILLCELL_X2 FILLER_75_694 ();
 FILLCELL_X2 FILLER_75_703 ();
 FILLCELL_X4 FILLER_75_712 ();
 FILLCELL_X2 FILLER_75_720 ();
 FILLCELL_X1 FILLER_75_722 ();
 FILLCELL_X4 FILLER_75_734 ();
 FILLCELL_X1 FILLER_75_742 ();
 FILLCELL_X1 FILLER_75_747 ();
 FILLCELL_X2 FILLER_75_756 ();
 FILLCELL_X1 FILLER_75_763 ();
 FILLCELL_X8 FILLER_75_771 ();
 FILLCELL_X1 FILLER_75_793 ();
 FILLCELL_X4 FILLER_75_808 ();
 FILLCELL_X2 FILLER_75_812 ();
 FILLCELL_X4 FILLER_75_821 ();
 FILLCELL_X1 FILLER_75_825 ();
 FILLCELL_X2 FILLER_75_875 ();
 FILLCELL_X2 FILLER_75_879 ();
 FILLCELL_X1 FILLER_75_885 ();
 FILLCELL_X2 FILLER_75_903 ();
 FILLCELL_X8 FILLER_75_917 ();
 FILLCELL_X4 FILLER_75_925 ();
 FILLCELL_X2 FILLER_75_929 ();
 FILLCELL_X1 FILLER_75_954 ();
 FILLCELL_X4 FILLER_75_960 ();
 FILLCELL_X2 FILLER_75_964 ();
 FILLCELL_X4 FILLER_75_973 ();
 FILLCELL_X16 FILLER_75_981 ();
 FILLCELL_X1 FILLER_75_997 ();
 FILLCELL_X1 FILLER_75_1003 ();
 FILLCELL_X1 FILLER_75_1008 ();
 FILLCELL_X1 FILLER_75_1013 ();
 FILLCELL_X2 FILLER_75_1020 ();
 FILLCELL_X4 FILLER_75_1028 ();
 FILLCELL_X4 FILLER_75_1060 ();
 FILLCELL_X2 FILLER_75_1064 ();
 FILLCELL_X4 FILLER_75_1072 ();
 FILLCELL_X2 FILLER_75_1082 ();
 FILLCELL_X1 FILLER_75_1084 ();
 FILLCELL_X2 FILLER_75_1113 ();
 FILLCELL_X1 FILLER_75_1115 ();
 FILLCELL_X2 FILLER_75_1118 ();
 FILLCELL_X4 FILLER_75_1123 ();
 FILLCELL_X1 FILLER_75_1127 ();
 FILLCELL_X1 FILLER_75_1135 ();
 FILLCELL_X4 FILLER_75_1168 ();
 FILLCELL_X1 FILLER_75_1172 ();
 FILLCELL_X2 FILLER_75_1193 ();
 FILLCELL_X1 FILLER_75_1236 ();
 FILLCELL_X4 FILLER_75_1249 ();
 FILLCELL_X2 FILLER_75_1253 ();
 FILLCELL_X2 FILLER_76_35 ();
 FILLCELL_X8 FILLER_76_44 ();
 FILLCELL_X8 FILLER_76_59 ();
 FILLCELL_X4 FILLER_76_67 ();
 FILLCELL_X2 FILLER_76_71 ();
 FILLCELL_X1 FILLER_76_73 ();
 FILLCELL_X16 FILLER_76_81 ();
 FILLCELL_X8 FILLER_76_97 ();
 FILLCELL_X4 FILLER_76_105 ();
 FILLCELL_X2 FILLER_76_109 ();
 FILLCELL_X2 FILLER_76_126 ();
 FILLCELL_X1 FILLER_76_128 ();
 FILLCELL_X16 FILLER_76_143 ();
 FILLCELL_X2 FILLER_76_159 ();
 FILLCELL_X1 FILLER_76_168 ();
 FILLCELL_X2 FILLER_76_189 ();
 FILLCELL_X2 FILLER_76_211 ();
 FILLCELL_X2 FILLER_76_217 ();
 FILLCELL_X4 FILLER_76_253 ();
 FILLCELL_X2 FILLER_76_257 ();
 FILLCELL_X1 FILLER_76_259 ();
 FILLCELL_X4 FILLER_76_287 ();
 FILLCELL_X1 FILLER_76_291 ();
 FILLCELL_X4 FILLER_76_296 ();
 FILLCELL_X2 FILLER_76_300 ();
 FILLCELL_X4 FILLER_76_305 ();
 FILLCELL_X2 FILLER_76_309 ();
 FILLCELL_X4 FILLER_76_323 ();
 FILLCELL_X2 FILLER_76_327 ();
 FILLCELL_X1 FILLER_76_329 ();
 FILLCELL_X8 FILLER_76_333 ();
 FILLCELL_X4 FILLER_76_341 ();
 FILLCELL_X2 FILLER_76_366 ();
 FILLCELL_X1 FILLER_76_368 ();
 FILLCELL_X4 FILLER_76_392 ();
 FILLCELL_X2 FILLER_76_396 ();
 FILLCELL_X4 FILLER_76_405 ();
 FILLCELL_X2 FILLER_76_409 ();
 FILLCELL_X2 FILLER_76_423 ();
 FILLCELL_X1 FILLER_76_445 ();
 FILLCELL_X1 FILLER_76_453 ();
 FILLCELL_X2 FILLER_76_458 ();
 FILLCELL_X4 FILLER_76_469 ();
 FILLCELL_X2 FILLER_76_473 ();
 FILLCELL_X1 FILLER_76_475 ();
 FILLCELL_X2 FILLER_76_487 ();
 FILLCELL_X2 FILLER_76_509 ();
 FILLCELL_X4 FILLER_76_530 ();
 FILLCELL_X4 FILLER_76_541 ();
 FILLCELL_X1 FILLER_76_545 ();
 FILLCELL_X4 FILLER_76_582 ();
 FILLCELL_X1 FILLER_76_586 ();
 FILLCELL_X4 FILLER_76_610 ();
 FILLCELL_X1 FILLER_76_637 ();
 FILLCELL_X1 FILLER_76_642 ();
 FILLCELL_X1 FILLER_76_653 ();
 FILLCELL_X8 FILLER_76_672 ();
 FILLCELL_X1 FILLER_76_680 ();
 FILLCELL_X2 FILLER_76_697 ();
 FILLCELL_X1 FILLER_76_699 ();
 FILLCELL_X2 FILLER_76_705 ();
 FILLCELL_X1 FILLER_76_707 ();
 FILLCELL_X4 FILLER_76_719 ();
 FILLCELL_X2 FILLER_76_723 ();
 FILLCELL_X1 FILLER_76_725 ();
 FILLCELL_X4 FILLER_76_731 ();
 FILLCELL_X2 FILLER_76_735 ();
 FILLCELL_X4 FILLER_76_751 ();
 FILLCELL_X2 FILLER_76_755 ();
 FILLCELL_X8 FILLER_76_786 ();
 FILLCELL_X2 FILLER_76_794 ();
 FILLCELL_X2 FILLER_76_801 ();
 FILLCELL_X4 FILLER_76_806 ();
 FILLCELL_X2 FILLER_76_810 ();
 FILLCELL_X4 FILLER_76_819 ();
 FILLCELL_X2 FILLER_76_823 ();
 FILLCELL_X4 FILLER_76_835 ();
 FILLCELL_X4 FILLER_76_847 ();
 FILLCELL_X2 FILLER_76_851 ();
 FILLCELL_X1 FILLER_76_860 ();
 FILLCELL_X4 FILLER_76_882 ();
 FILLCELL_X2 FILLER_76_886 ();
 FILLCELL_X1 FILLER_76_888 ();
 FILLCELL_X8 FILLER_76_893 ();
 FILLCELL_X1 FILLER_76_901 ();
 FILLCELL_X4 FILLER_76_918 ();
 FILLCELL_X1 FILLER_76_922 ();
 FILLCELL_X2 FILLER_76_944 ();
 FILLCELL_X8 FILLER_76_986 ();
 FILLCELL_X4 FILLER_76_994 ();
 FILLCELL_X2 FILLER_76_998 ();
 FILLCELL_X1 FILLER_76_1000 ();
 FILLCELL_X8 FILLER_76_1022 ();
 FILLCELL_X1 FILLER_76_1030 ();
 FILLCELL_X2 FILLER_76_1062 ();
 FILLCELL_X1 FILLER_76_1064 ();
 FILLCELL_X16 FILLER_76_1083 ();
 FILLCELL_X1 FILLER_76_1103 ();
 FILLCELL_X4 FILLER_76_1108 ();
 FILLCELL_X2 FILLER_76_1112 ();
 FILLCELL_X1 FILLER_76_1140 ();
 FILLCELL_X1 FILLER_76_1158 ();
 FILLCELL_X2 FILLER_76_1169 ();
 FILLCELL_X4 FILLER_76_1176 ();
 FILLCELL_X2 FILLER_76_1180 ();
 FILLCELL_X4 FILLER_76_1195 ();
 FILLCELL_X2 FILLER_76_1199 ();
 FILLCELL_X1 FILLER_76_1201 ();
 FILLCELL_X4 FILLER_76_1212 ();
 FILLCELL_X2 FILLER_76_1216 ();
 FILLCELL_X4 FILLER_76_1222 ();
 FILLCELL_X16 FILLER_76_1234 ();
 FILLCELL_X1 FILLER_76_1250 ();
 FILLCELL_X2 FILLER_77_1 ();
 FILLCELL_X4 FILLER_77_8 ();
 FILLCELL_X2 FILLER_77_12 ();
 FILLCELL_X1 FILLER_77_34 ();
 FILLCELL_X2 FILLER_77_42 ();
 FILLCELL_X1 FILLER_77_44 ();
 FILLCELL_X1 FILLER_77_55 ();
 FILLCELL_X2 FILLER_77_63 ();
 FILLCELL_X1 FILLER_77_65 ();
 FILLCELL_X8 FILLER_77_73 ();
 FILLCELL_X4 FILLER_77_81 ();
 FILLCELL_X1 FILLER_77_85 ();
 FILLCELL_X4 FILLER_77_93 ();
 FILLCELL_X2 FILLER_77_97 ();
 FILLCELL_X16 FILLER_77_174 ();
 FILLCELL_X4 FILLER_77_190 ();
 FILLCELL_X2 FILLER_77_196 ();
 FILLCELL_X2 FILLER_77_226 ();
 FILLCELL_X2 FILLER_77_263 ();
 FILLCELL_X1 FILLER_77_265 ();
 FILLCELL_X4 FILLER_77_277 ();
 FILLCELL_X2 FILLER_77_281 ();
 FILLCELL_X1 FILLER_77_286 ();
 FILLCELL_X4 FILLER_77_330 ();
 FILLCELL_X2 FILLER_77_334 ();
 FILLCELL_X1 FILLER_77_389 ();
 FILLCELL_X4 FILLER_77_413 ();
 FILLCELL_X2 FILLER_77_417 ();
 FILLCELL_X1 FILLER_77_493 ();
 FILLCELL_X8 FILLER_77_510 ();
 FILLCELL_X8 FILLER_77_525 ();
 FILLCELL_X4 FILLER_77_533 ();
 FILLCELL_X2 FILLER_77_537 ();
 FILLCELL_X1 FILLER_77_559 ();
 FILLCELL_X4 FILLER_77_609 ();
 FILLCELL_X2 FILLER_77_613 ();
 FILLCELL_X1 FILLER_77_615 ();
 FILLCELL_X1 FILLER_77_659 ();
 FILLCELL_X2 FILLER_77_662 ();
 FILLCELL_X1 FILLER_77_664 ();
 FILLCELL_X16 FILLER_77_682 ();
 FILLCELL_X4 FILLER_77_698 ();
 FILLCELL_X8 FILLER_77_714 ();
 FILLCELL_X2 FILLER_77_722 ();
 FILLCELL_X1 FILLER_77_724 ();
 FILLCELL_X1 FILLER_77_732 ();
 FILLCELL_X2 FILLER_77_736 ();
 FILLCELL_X2 FILLER_77_744 ();
 FILLCELL_X4 FILLER_77_753 ();
 FILLCELL_X2 FILLER_77_774 ();
 FILLCELL_X4 FILLER_77_785 ();
 FILLCELL_X2 FILLER_77_810 ();
 FILLCELL_X1 FILLER_77_812 ();
 FILLCELL_X4 FILLER_77_820 ();
 FILLCELL_X2 FILLER_77_824 ();
 FILLCELL_X1 FILLER_77_826 ();
 FILLCELL_X2 FILLER_77_840 ();
 FILLCELL_X2 FILLER_77_849 ();
 FILLCELL_X1 FILLER_77_851 ();
 FILLCELL_X4 FILLER_77_902 ();
 FILLCELL_X16 FILLER_77_913 ();
 FILLCELL_X2 FILLER_77_936 ();
 FILLCELL_X4 FILLER_77_945 ();
 FILLCELL_X4 FILLER_77_956 ();
 FILLCELL_X4 FILLER_77_962 ();
 FILLCELL_X2 FILLER_77_966 ();
 FILLCELL_X4 FILLER_77_977 ();
 FILLCELL_X1 FILLER_77_981 ();
 FILLCELL_X8 FILLER_77_999 ();
 FILLCELL_X2 FILLER_77_1018 ();
 FILLCELL_X4 FILLER_77_1051 ();
 FILLCELL_X1 FILLER_77_1055 ();
 FILLCELL_X1 FILLER_77_1076 ();
 FILLCELL_X4 FILLER_77_1091 ();
 FILLCELL_X1 FILLER_77_1095 ();
 FILLCELL_X4 FILLER_77_1110 ();
 FILLCELL_X1 FILLER_77_1114 ();
 FILLCELL_X16 FILLER_77_1122 ();
 FILLCELL_X2 FILLER_77_1138 ();
 FILLCELL_X1 FILLER_77_1140 ();
 FILLCELL_X4 FILLER_77_1155 ();
 FILLCELL_X1 FILLER_77_1162 ();
 FILLCELL_X1 FILLER_77_1185 ();
 FILLCELL_X1 FILLER_77_1201 ();
 FILLCELL_X4 FILLER_77_1207 ();
 FILLCELL_X1 FILLER_77_1211 ();
 FILLCELL_X2 FILLER_77_1215 ();
 FILLCELL_X1 FILLER_77_1217 ();
 FILLCELL_X2 FILLER_77_1243 ();
 FILLCELL_X1 FILLER_77_1245 ();
 FILLCELL_X1 FILLER_77_1249 ();
 FILLCELL_X2 FILLER_77_1253 ();
 FILLCELL_X8 FILLER_78_1 ();
 FILLCELL_X4 FILLER_78_9 ();
 FILLCELL_X2 FILLER_78_13 ();
 FILLCELL_X2 FILLER_78_22 ();
 FILLCELL_X4 FILLER_78_38 ();
 FILLCELL_X2 FILLER_78_42 ();
 FILLCELL_X4 FILLER_78_104 ();
 FILLCELL_X2 FILLER_78_108 ();
 FILLCELL_X1 FILLER_78_110 ();
 FILLCELL_X4 FILLER_78_118 ();
 FILLCELL_X1 FILLER_78_122 ();
 FILLCELL_X1 FILLER_78_135 ();
 FILLCELL_X8 FILLER_78_143 ();
 FILLCELL_X1 FILLER_78_151 ();
 FILLCELL_X2 FILLER_78_155 ();
 FILLCELL_X8 FILLER_78_164 ();
 FILLCELL_X2 FILLER_78_176 ();
 FILLCELL_X1 FILLER_78_178 ();
 FILLCELL_X2 FILLER_78_201 ();
 FILLCELL_X1 FILLER_78_206 ();
 FILLCELL_X4 FILLER_78_215 ();
 FILLCELL_X2 FILLER_78_219 ();
 FILLCELL_X4 FILLER_78_225 ();
 FILLCELL_X2 FILLER_78_229 ();
 FILLCELL_X32 FILLER_78_234 ();
 FILLCELL_X2 FILLER_78_270 ();
 FILLCELL_X1 FILLER_78_272 ();
 FILLCELL_X2 FILLER_78_276 ();
 FILLCELL_X4 FILLER_78_285 ();
 FILLCELL_X2 FILLER_78_293 ();
 FILLCELL_X8 FILLER_78_302 ();
 FILLCELL_X1 FILLER_78_310 ();
 FILLCELL_X1 FILLER_78_333 ();
 FILLCELL_X4 FILLER_78_354 ();
 FILLCELL_X1 FILLER_78_358 ();
 FILLCELL_X2 FILLER_78_373 ();
 FILLCELL_X4 FILLER_78_388 ();
 FILLCELL_X2 FILLER_78_396 ();
 FILLCELL_X2 FILLER_78_409 ();
 FILLCELL_X2 FILLER_78_438 ();
 FILLCELL_X1 FILLER_78_440 ();
 FILLCELL_X4 FILLER_78_448 ();
 FILLCELL_X8 FILLER_78_459 ();
 FILLCELL_X2 FILLER_78_467 ();
 FILLCELL_X1 FILLER_78_469 ();
 FILLCELL_X4 FILLER_78_473 ();
 FILLCELL_X2 FILLER_78_477 ();
 FILLCELL_X1 FILLER_78_479 ();
 FILLCELL_X4 FILLER_78_484 ();
 FILLCELL_X2 FILLER_78_488 ();
 FILLCELL_X4 FILLER_78_525 ();
 FILLCELL_X2 FILLER_78_529 ();
 FILLCELL_X1 FILLER_78_531 ();
 FILLCELL_X8 FILLER_78_544 ();
 FILLCELL_X1 FILLER_78_552 ();
 FILLCELL_X8 FILLER_78_572 ();
 FILLCELL_X4 FILLER_78_580 ();
 FILLCELL_X2 FILLER_78_584 ();
 FILLCELL_X1 FILLER_78_586 ();
 FILLCELL_X16 FILLER_78_594 ();
 FILLCELL_X2 FILLER_78_610 ();
 FILLCELL_X2 FILLER_78_619 ();
 FILLCELL_X1 FILLER_78_621 ();
 FILLCELL_X4 FILLER_78_624 ();
 FILLCELL_X2 FILLER_78_628 ();
 FILLCELL_X1 FILLER_78_630 ();
 FILLCELL_X8 FILLER_78_632 ();
 FILLCELL_X1 FILLER_78_640 ();
 FILLCELL_X2 FILLER_78_667 ();
 FILLCELL_X8 FILLER_78_682 ();
 FILLCELL_X4 FILLER_78_690 ();
 FILLCELL_X1 FILLER_78_694 ();
 FILLCELL_X4 FILLER_78_717 ();
 FILLCELL_X2 FILLER_78_721 ();
 FILLCELL_X1 FILLER_78_743 ();
 FILLCELL_X1 FILLER_78_759 ();
 FILLCELL_X2 FILLER_78_765 ();
 FILLCELL_X1 FILLER_78_771 ();
 FILLCELL_X2 FILLER_78_783 ();
 FILLCELL_X4 FILLER_78_792 ();
 FILLCELL_X1 FILLER_78_807 ();
 FILLCELL_X2 FILLER_78_840 ();
 FILLCELL_X1 FILLER_78_842 ();
 FILLCELL_X16 FILLER_78_846 ();
 FILLCELL_X4 FILLER_78_862 ();
 FILLCELL_X32 FILLER_78_871 ();
 FILLCELL_X4 FILLER_78_903 ();
 FILLCELL_X1 FILLER_78_907 ();
 FILLCELL_X2 FILLER_78_970 ();
 FILLCELL_X2 FILLER_78_994 ();
 FILLCELL_X1 FILLER_78_1013 ();
 FILLCELL_X8 FILLER_78_1017 ();
 FILLCELL_X4 FILLER_78_1025 ();
 FILLCELL_X1 FILLER_78_1029 ();
 FILLCELL_X2 FILLER_78_1044 ();
 FILLCELL_X1 FILLER_78_1046 ();
 FILLCELL_X8 FILLER_78_1054 ();
 FILLCELL_X8 FILLER_78_1085 ();
 FILLCELL_X4 FILLER_78_1093 ();
 FILLCELL_X1 FILLER_78_1097 ();
 FILLCELL_X4 FILLER_78_1111 ();
 FILLCELL_X2 FILLER_78_1115 ();
 FILLCELL_X1 FILLER_78_1117 ();
 FILLCELL_X4 FILLER_78_1125 ();
 FILLCELL_X2 FILLER_78_1129 ();
 FILLCELL_X1 FILLER_78_1131 ();
 FILLCELL_X2 FILLER_78_1139 ();
 FILLCELL_X1 FILLER_78_1145 ();
 FILLCELL_X1 FILLER_78_1151 ();
 FILLCELL_X1 FILLER_78_1166 ();
 FILLCELL_X1 FILLER_78_1169 ();
 FILLCELL_X2 FILLER_78_1176 ();
 FILLCELL_X2 FILLER_78_1199 ();
 FILLCELL_X1 FILLER_78_1211 ();
 FILLCELL_X1 FILLER_78_1217 ();
 FILLCELL_X2 FILLER_78_1224 ();
 FILLCELL_X1 FILLER_79_28 ();
 FILLCELL_X2 FILLER_79_43 ();
 FILLCELL_X1 FILLER_79_45 ();
 FILLCELL_X1 FILLER_79_58 ();
 FILLCELL_X2 FILLER_79_66 ();
 FILLCELL_X2 FILLER_79_75 ();
 FILLCELL_X1 FILLER_79_77 ();
 FILLCELL_X1 FILLER_79_85 ();
 FILLCELL_X2 FILLER_79_93 ();
 FILLCELL_X1 FILLER_79_95 ();
 FILLCELL_X2 FILLER_79_180 ();
 FILLCELL_X4 FILLER_79_185 ();
 FILLCELL_X1 FILLER_79_200 ();
 FILLCELL_X1 FILLER_79_205 ();
 FILLCELL_X4 FILLER_79_210 ();
 FILLCELL_X1 FILLER_79_214 ();
 FILLCELL_X4 FILLER_79_235 ();
 FILLCELL_X2 FILLER_79_253 ();
 FILLCELL_X1 FILLER_79_287 ();
 FILLCELL_X2 FILLER_79_304 ();
 FILLCELL_X1 FILLER_79_306 ();
 FILLCELL_X8 FILLER_79_310 ();
 FILLCELL_X1 FILLER_79_318 ();
 FILLCELL_X8 FILLER_79_330 ();
 FILLCELL_X1 FILLER_79_338 ();
 FILLCELL_X4 FILLER_79_365 ();
 FILLCELL_X1 FILLER_79_369 ();
 FILLCELL_X8 FILLER_79_405 ();
 FILLCELL_X2 FILLER_79_413 ();
 FILLCELL_X1 FILLER_79_415 ();
 FILLCELL_X1 FILLER_79_429 ();
 FILLCELL_X2 FILLER_79_470 ();
 FILLCELL_X8 FILLER_79_479 ();
 FILLCELL_X1 FILLER_79_487 ();
 FILLCELL_X8 FILLER_79_493 ();
 FILLCELL_X8 FILLER_79_511 ();
 FILLCELL_X2 FILLER_79_519 ();
 FILLCELL_X1 FILLER_79_521 ();
 FILLCELL_X1 FILLER_79_555 ();
 FILLCELL_X4 FILLER_79_570 ();
 FILLCELL_X1 FILLER_79_574 ();
 FILLCELL_X8 FILLER_79_582 ();
 FILLCELL_X1 FILLER_79_590 ();
 FILLCELL_X8 FILLER_79_605 ();
 FILLCELL_X4 FILLER_79_613 ();
 FILLCELL_X2 FILLER_79_617 ();
 FILLCELL_X1 FILLER_79_619 ();
 FILLCELL_X2 FILLER_79_630 ();
 FILLCELL_X2 FILLER_79_646 ();
 FILLCELL_X8 FILLER_79_673 ();
 FILLCELL_X4 FILLER_79_681 ();
 FILLCELL_X8 FILLER_79_702 ();
 FILLCELL_X1 FILLER_79_710 ();
 FILLCELL_X4 FILLER_79_731 ();
 FILLCELL_X2 FILLER_79_735 ();
 FILLCELL_X1 FILLER_79_737 ();
 FILLCELL_X2 FILLER_79_750 ();
 FILLCELL_X1 FILLER_79_752 ();
 FILLCELL_X4 FILLER_79_758 ();
 FILLCELL_X2 FILLER_79_762 ();
 FILLCELL_X2 FILLER_79_781 ();
 FILLCELL_X1 FILLER_79_783 ();
 FILLCELL_X4 FILLER_79_791 ();
 FILLCELL_X2 FILLER_79_795 ();
 FILLCELL_X8 FILLER_79_811 ();
 FILLCELL_X4 FILLER_79_826 ();
 FILLCELL_X2 FILLER_79_830 ();
 FILLCELL_X1 FILLER_79_832 ();
 FILLCELL_X16 FILLER_79_842 ();
 FILLCELL_X4 FILLER_79_858 ();
 FILLCELL_X2 FILLER_79_862 ();
 FILLCELL_X1 FILLER_79_864 ();
 FILLCELL_X16 FILLER_79_885 ();
 FILLCELL_X2 FILLER_79_901 ();
 FILLCELL_X1 FILLER_79_903 ();
 FILLCELL_X4 FILLER_79_909 ();
 FILLCELL_X2 FILLER_79_920 ();
 FILLCELL_X2 FILLER_79_931 ();
 FILLCELL_X1 FILLER_79_933 ();
 FILLCELL_X2 FILLER_79_941 ();
 FILLCELL_X1 FILLER_79_943 ();
 FILLCELL_X2 FILLER_79_958 ();
 FILLCELL_X8 FILLER_79_963 ();
 FILLCELL_X2 FILLER_79_971 ();
 FILLCELL_X1 FILLER_79_973 ();
 FILLCELL_X2 FILLER_79_979 ();
 FILLCELL_X8 FILLER_79_992 ();
 FILLCELL_X2 FILLER_79_1000 ();
 FILLCELL_X1 FILLER_79_1002 ();
 FILLCELL_X4 FILLER_79_1030 ();
 FILLCELL_X1 FILLER_79_1034 ();
 FILLCELL_X1 FILLER_79_1042 ();
 FILLCELL_X2 FILLER_79_1049 ();
 FILLCELL_X1 FILLER_79_1051 ();
 FILLCELL_X2 FILLER_79_1059 ();
 FILLCELL_X1 FILLER_79_1061 ();
 FILLCELL_X4 FILLER_79_1076 ();
 FILLCELL_X1 FILLER_79_1080 ();
 FILLCELL_X2 FILLER_79_1095 ();
 FILLCELL_X2 FILLER_79_1103 ();
 FILLCELL_X1 FILLER_79_1105 ();
 FILLCELL_X1 FILLER_79_1110 ();
 FILLCELL_X2 FILLER_79_1128 ();
 FILLCELL_X1 FILLER_79_1130 ();
 FILLCELL_X1 FILLER_79_1140 ();
 FILLCELL_X2 FILLER_79_1158 ();
 FILLCELL_X1 FILLER_79_1160 ();
 FILLCELL_X2 FILLER_79_1167 ();
 FILLCELL_X1 FILLER_79_1169 ();
 FILLCELL_X16 FILLER_79_1178 ();
 FILLCELL_X2 FILLER_79_1194 ();
 FILLCELL_X2 FILLER_79_1199 ();
 FILLCELL_X2 FILLER_79_1206 ();
 FILLCELL_X1 FILLER_79_1213 ();
 FILLCELL_X1 FILLER_79_1220 ();
 FILLCELL_X4 FILLER_79_1238 ();
 FILLCELL_X2 FILLER_79_1242 ();
 FILLCELL_X1 FILLER_79_1244 ();
 FILLCELL_X2 FILLER_79_1248 ();
 FILLCELL_X1 FILLER_79_1254 ();
 FILLCELL_X8 FILLER_80_1 ();
 FILLCELL_X4 FILLER_80_9 ();
 FILLCELL_X2 FILLER_80_13 ();
 FILLCELL_X8 FILLER_80_42 ();
 FILLCELL_X1 FILLER_80_77 ();
 FILLCELL_X1 FILLER_80_85 ();
 FILLCELL_X2 FILLER_80_93 ();
 FILLCELL_X1 FILLER_80_115 ();
 FILLCELL_X8 FILLER_80_123 ();
 FILLCELL_X16 FILLER_80_138 ();
 FILLCELL_X2 FILLER_80_154 ();
 FILLCELL_X1 FILLER_80_156 ();
 FILLCELL_X4 FILLER_80_164 ();
 FILLCELL_X2 FILLER_80_168 ();
 FILLCELL_X1 FILLER_80_170 ();
 FILLCELL_X1 FILLER_80_181 ();
 FILLCELL_X1 FILLER_80_185 ();
 FILLCELL_X4 FILLER_80_203 ();
 FILLCELL_X1 FILLER_80_207 ();
 FILLCELL_X4 FILLER_80_218 ();
 FILLCELL_X2 FILLER_80_222 ();
 FILLCELL_X1 FILLER_80_224 ();
 FILLCELL_X1 FILLER_80_232 ();
 FILLCELL_X4 FILLER_80_256 ();
 FILLCELL_X8 FILLER_80_276 ();
 FILLCELL_X2 FILLER_80_287 ();
 FILLCELL_X1 FILLER_80_293 ();
 FILLCELL_X1 FILLER_80_311 ();
 FILLCELL_X1 FILLER_80_316 ();
 FILLCELL_X8 FILLER_80_327 ();
 FILLCELL_X4 FILLER_80_369 ();
 FILLCELL_X1 FILLER_80_373 ();
 FILLCELL_X2 FILLER_80_431 ();
 FILLCELL_X2 FILLER_80_436 ();
 FILLCELL_X1 FILLER_80_438 ();
 FILLCELL_X2 FILLER_80_442 ();
 FILLCELL_X1 FILLER_80_444 ();
 FILLCELL_X1 FILLER_80_454 ();
 FILLCELL_X2 FILLER_80_476 ();
 FILLCELL_X2 FILLER_80_498 ();
 FILLCELL_X2 FILLER_80_509 ();
 FILLCELL_X1 FILLER_80_511 ();
 FILLCELL_X4 FILLER_80_519 ();
 FILLCELL_X2 FILLER_80_523 ();
 FILLCELL_X1 FILLER_80_525 ();
 FILLCELL_X8 FILLER_80_546 ();
 FILLCELL_X4 FILLER_80_561 ();
 FILLCELL_X2 FILLER_80_565 ();
 FILLCELL_X1 FILLER_80_567 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X4 FILLER_80_632 ();
 FILLCELL_X1 FILLER_80_636 ();
 FILLCELL_X4 FILLER_80_651 ();
 FILLCELL_X2 FILLER_80_655 ();
 FILLCELL_X1 FILLER_80_657 ();
 FILLCELL_X4 FILLER_80_663 ();
 FILLCELL_X1 FILLER_80_667 ();
 FILLCELL_X4 FILLER_80_690 ();
 FILLCELL_X1 FILLER_80_694 ();
 FILLCELL_X1 FILLER_80_711 ();
 FILLCELL_X1 FILLER_80_715 ();
 FILLCELL_X2 FILLER_80_723 ();
 FILLCELL_X8 FILLER_80_754 ();
 FILLCELL_X4 FILLER_80_762 ();
 FILLCELL_X2 FILLER_80_766 ();
 FILLCELL_X2 FILLER_80_781 ();
 FILLCELL_X1 FILLER_80_783 ();
 FILLCELL_X2 FILLER_80_795 ();
 FILLCELL_X1 FILLER_80_797 ();
 FILLCELL_X8 FILLER_80_807 ();
 FILLCELL_X2 FILLER_80_815 ();
 FILLCELL_X8 FILLER_80_834 ();
 FILLCELL_X4 FILLER_80_842 ();
 FILLCELL_X2 FILLER_80_846 ();
 FILLCELL_X1 FILLER_80_848 ();
 FILLCELL_X16 FILLER_80_873 ();
 FILLCELL_X4 FILLER_80_889 ();
 FILLCELL_X2 FILLER_80_893 ();
 FILLCELL_X4 FILLER_80_902 ();
 FILLCELL_X2 FILLER_80_906 ();
 FILLCELL_X2 FILLER_80_919 ();
 FILLCELL_X1 FILLER_80_921 ();
 FILLCELL_X1 FILLER_80_940 ();
 FILLCELL_X1 FILLER_80_982 ();
 FILLCELL_X8 FILLER_80_1006 ();
 FILLCELL_X2 FILLER_80_1014 ();
 FILLCELL_X1 FILLER_80_1016 ();
 FILLCELL_X1 FILLER_80_1020 ();
 FILLCELL_X1 FILLER_80_1054 ();
 FILLCELL_X1 FILLER_80_1076 ();
 FILLCELL_X2 FILLER_80_1082 ();
 FILLCELL_X2 FILLER_80_1090 ();
 FILLCELL_X2 FILLER_80_1099 ();
 FILLCELL_X2 FILLER_80_1141 ();
 FILLCELL_X4 FILLER_80_1147 ();
 FILLCELL_X1 FILLER_80_1163 ();
 FILLCELL_X1 FILLER_80_1208 ();
 FILLCELL_X1 FILLER_80_1215 ();
 FILLCELL_X1 FILLER_80_1220 ();
 FILLCELL_X4 FILLER_80_1225 ();
 FILLCELL_X4 FILLER_80_1232 ();
 FILLCELL_X1 FILLER_80_1236 ();
 FILLCELL_X4 FILLER_80_1240 ();
 FILLCELL_X4 FILLER_80_1248 ();
 FILLCELL_X2 FILLER_80_1252 ();
 FILLCELL_X1 FILLER_80_1254 ();
 FILLCELL_X1 FILLER_81_1 ();
 FILLCELL_X4 FILLER_81_22 ();
 FILLCELL_X2 FILLER_81_26 ();
 FILLCELL_X4 FILLER_81_48 ();
 FILLCELL_X1 FILLER_81_52 ();
 FILLCELL_X8 FILLER_81_67 ();
 FILLCELL_X4 FILLER_81_75 ();
 FILLCELL_X2 FILLER_81_79 ();
 FILLCELL_X16 FILLER_81_88 ();
 FILLCELL_X4 FILLER_81_158 ();
 FILLCELL_X1 FILLER_81_169 ();
 FILLCELL_X4 FILLER_81_180 ();
 FILLCELL_X2 FILLER_81_188 ();
 FILLCELL_X8 FILLER_81_194 ();
 FILLCELL_X1 FILLER_81_202 ();
 FILLCELL_X2 FILLER_81_217 ();
 FILLCELL_X1 FILLER_81_219 ();
 FILLCELL_X2 FILLER_81_227 ();
 FILLCELL_X1 FILLER_81_249 ();
 FILLCELL_X2 FILLER_81_257 ();
 FILLCELL_X1 FILLER_81_263 ();
 FILLCELL_X4 FILLER_81_267 ();
 FILLCELL_X2 FILLER_81_275 ();
 FILLCELL_X1 FILLER_81_277 ();
 FILLCELL_X2 FILLER_81_281 ();
 FILLCELL_X2 FILLER_81_303 ();
 FILLCELL_X4 FILLER_81_339 ();
 FILLCELL_X1 FILLER_81_343 ();
 FILLCELL_X1 FILLER_81_349 ();
 FILLCELL_X4 FILLER_81_397 ();
 FILLCELL_X1 FILLER_81_401 ();
 FILLCELL_X16 FILLER_81_431 ();
 FILLCELL_X1 FILLER_81_447 ();
 FILLCELL_X2 FILLER_81_460 ();
 FILLCELL_X8 FILLER_81_469 ();
 FILLCELL_X4 FILLER_81_503 ();
 FILLCELL_X2 FILLER_81_507 ();
 FILLCELL_X16 FILLER_81_518 ();
 FILLCELL_X8 FILLER_81_534 ();
 FILLCELL_X1 FILLER_81_542 ();
 FILLCELL_X1 FILLER_81_547 ();
 FILLCELL_X1 FILLER_81_568 ();
 FILLCELL_X4 FILLER_81_603 ();
 FILLCELL_X2 FILLER_81_607 ();
 FILLCELL_X1 FILLER_81_609 ();
 FILLCELL_X1 FILLER_81_624 ();
 FILLCELL_X8 FILLER_81_638 ();
 FILLCELL_X8 FILLER_81_653 ();
 FILLCELL_X4 FILLER_81_661 ();
 FILLCELL_X16 FILLER_81_674 ();
 FILLCELL_X8 FILLER_81_690 ();
 FILLCELL_X2 FILLER_81_698 ();
 FILLCELL_X2 FILLER_81_707 ();
 FILLCELL_X2 FILLER_81_730 ();
 FILLCELL_X1 FILLER_81_759 ();
 FILLCELL_X8 FILLER_81_764 ();
 FILLCELL_X4 FILLER_81_772 ();
 FILLCELL_X2 FILLER_81_794 ();
 FILLCELL_X1 FILLER_81_796 ();
 FILLCELL_X4 FILLER_81_801 ();
 FILLCELL_X4 FILLER_81_815 ();
 FILLCELL_X4 FILLER_81_822 ();
 FILLCELL_X1 FILLER_81_826 ();
 FILLCELL_X1 FILLER_81_842 ();
 FILLCELL_X2 FILLER_81_860 ();
 FILLCELL_X1 FILLER_81_865 ();
 FILLCELL_X2 FILLER_81_876 ();
 FILLCELL_X1 FILLER_81_914 ();
 FILLCELL_X1 FILLER_81_933 ();
 FILLCELL_X16 FILLER_81_944 ();
 FILLCELL_X8 FILLER_81_960 ();
 FILLCELL_X2 FILLER_81_968 ();
 FILLCELL_X16 FILLER_81_992 ();
 FILLCELL_X8 FILLER_81_1008 ();
 FILLCELL_X2 FILLER_81_1016 ();
 FILLCELL_X1 FILLER_81_1018 ();
 FILLCELL_X1 FILLER_81_1022 ();
 FILLCELL_X2 FILLER_81_1026 ();
 FILLCELL_X8 FILLER_81_1031 ();
 FILLCELL_X4 FILLER_81_1039 ();
 FILLCELL_X2 FILLER_81_1043 ();
 FILLCELL_X1 FILLER_81_1045 ();
 FILLCELL_X16 FILLER_81_1056 ();
 FILLCELL_X4 FILLER_81_1072 ();
 FILLCELL_X2 FILLER_81_1076 ();
 FILLCELL_X1 FILLER_81_1078 ();
 FILLCELL_X1 FILLER_81_1094 ();
 FILLCELL_X8 FILLER_81_1114 ();
 FILLCELL_X2 FILLER_81_1122 ();
 FILLCELL_X1 FILLER_81_1124 ();
 FILLCELL_X16 FILLER_81_1134 ();
 FILLCELL_X2 FILLER_81_1150 ();
 FILLCELL_X1 FILLER_81_1156 ();
 FILLCELL_X8 FILLER_81_1166 ();
 FILLCELL_X2 FILLER_81_1174 ();
 FILLCELL_X1 FILLER_81_1176 ();
 FILLCELL_X4 FILLER_81_1190 ();
 FILLCELL_X2 FILLER_81_1194 ();
 FILLCELL_X4 FILLER_81_1203 ();
 FILLCELL_X8 FILLER_81_1215 ();
 FILLCELL_X2 FILLER_81_1223 ();
 FILLCELL_X1 FILLER_81_1225 ();
 FILLCELL_X4 FILLER_81_1247 ();
 FILLCELL_X1 FILLER_81_1251 ();
 FILLCELL_X8 FILLER_82_1 ();
 FILLCELL_X2 FILLER_82_9 ();
 FILLCELL_X8 FILLER_82_18 ();
 FILLCELL_X2 FILLER_82_26 ();
 FILLCELL_X1 FILLER_82_35 ();
 FILLCELL_X16 FILLER_82_70 ();
 FILLCELL_X1 FILLER_82_86 ();
 FILLCELL_X16 FILLER_82_121 ();
 FILLCELL_X8 FILLER_82_137 ();
 FILLCELL_X8 FILLER_82_152 ();
 FILLCELL_X2 FILLER_82_160 ();
 FILLCELL_X1 FILLER_82_162 ();
 FILLCELL_X2 FILLER_82_187 ();
 FILLCELL_X1 FILLER_82_189 ();
 FILLCELL_X8 FILLER_82_208 ();
 FILLCELL_X2 FILLER_82_216 ();
 FILLCELL_X1 FILLER_82_218 ();
 FILLCELL_X2 FILLER_82_229 ();
 FILLCELL_X4 FILLER_82_307 ();
 FILLCELL_X2 FILLER_82_311 ();
 FILLCELL_X2 FILLER_82_356 ();
 FILLCELL_X1 FILLER_82_379 ();
 FILLCELL_X4 FILLER_82_384 ();
 FILLCELL_X2 FILLER_82_399 ();
 FILLCELL_X4 FILLER_82_421 ();
 FILLCELL_X2 FILLER_82_425 ();
 FILLCELL_X1 FILLER_82_427 ();
 FILLCELL_X1 FILLER_82_432 ();
 FILLCELL_X1 FILLER_82_436 ();
 FILLCELL_X1 FILLER_82_464 ();
 FILLCELL_X4 FILLER_82_478 ();
 FILLCELL_X2 FILLER_82_482 ();
 FILLCELL_X8 FILLER_82_491 ();
 FILLCELL_X1 FILLER_82_499 ();
 FILLCELL_X1 FILLER_82_507 ();
 FILLCELL_X2 FILLER_82_535 ();
 FILLCELL_X2 FILLER_82_541 ();
 FILLCELL_X1 FILLER_82_543 ();
 FILLCELL_X2 FILLER_82_564 ();
 FILLCELL_X1 FILLER_82_566 ();
 FILLCELL_X32 FILLER_82_584 ();
 FILLCELL_X4 FILLER_82_616 ();
 FILLCELL_X2 FILLER_82_620 ();
 FILLCELL_X4 FILLER_82_632 ();
 FILLCELL_X1 FILLER_82_636 ();
 FILLCELL_X8 FILLER_82_673 ();
 FILLCELL_X1 FILLER_82_681 ();
 FILLCELL_X4 FILLER_82_689 ();
 FILLCELL_X2 FILLER_82_693 ();
 FILLCELL_X1 FILLER_82_695 ();
 FILLCELL_X1 FILLER_82_703 ();
 FILLCELL_X1 FILLER_82_719 ();
 FILLCELL_X4 FILLER_82_731 ();
 FILLCELL_X1 FILLER_82_735 ();
 FILLCELL_X2 FILLER_82_745 ();
 FILLCELL_X2 FILLER_82_751 ();
 FILLCELL_X1 FILLER_82_753 ();
 FILLCELL_X4 FILLER_82_765 ();
 FILLCELL_X2 FILLER_82_769 ();
 FILLCELL_X2 FILLER_82_778 ();
 FILLCELL_X2 FILLER_82_787 ();
 FILLCELL_X1 FILLER_82_789 ();
 FILLCELL_X1 FILLER_82_796 ();
 FILLCELL_X1 FILLER_82_808 ();
 FILLCELL_X4 FILLER_82_820 ();
 FILLCELL_X2 FILLER_82_824 ();
 FILLCELL_X1 FILLER_82_826 ();
 FILLCELL_X2 FILLER_82_838 ();
 FILLCELL_X4 FILLER_82_858 ();
 FILLCELL_X1 FILLER_82_862 ();
 FILLCELL_X2 FILLER_82_867 ();
 FILLCELL_X1 FILLER_82_869 ();
 FILLCELL_X2 FILLER_82_877 ();
 FILLCELL_X16 FILLER_82_889 ();
 FILLCELL_X8 FILLER_82_905 ();
 FILLCELL_X4 FILLER_82_913 ();
 FILLCELL_X1 FILLER_82_917 ();
 FILLCELL_X4 FILLER_82_924 ();
 FILLCELL_X1 FILLER_82_928 ();
 FILLCELL_X4 FILLER_82_946 ();
 FILLCELL_X2 FILLER_82_950 ();
 FILLCELL_X1 FILLER_82_952 ();
 FILLCELL_X8 FILLER_82_964 ();
 FILLCELL_X4 FILLER_82_972 ();
 FILLCELL_X1 FILLER_82_976 ();
 FILLCELL_X8 FILLER_82_997 ();
 FILLCELL_X2 FILLER_82_1005 ();
 FILLCELL_X2 FILLER_82_1012 ();
 FILLCELL_X1 FILLER_82_1014 ();
 FILLCELL_X2 FILLER_82_1018 ();
 FILLCELL_X4 FILLER_82_1044 ();
 FILLCELL_X8 FILLER_82_1065 ();
 FILLCELL_X2 FILLER_82_1095 ();
 FILLCELL_X1 FILLER_82_1097 ();
 FILLCELL_X2 FILLER_82_1115 ();
 FILLCELL_X1 FILLER_82_1117 ();
 FILLCELL_X2 FILLER_82_1125 ();
 FILLCELL_X1 FILLER_82_1127 ();
 FILLCELL_X4 FILLER_82_1135 ();
 FILLCELL_X1 FILLER_82_1139 ();
 FILLCELL_X1 FILLER_82_1145 ();
 FILLCELL_X8 FILLER_82_1186 ();
 FILLCELL_X4 FILLER_82_1194 ();
 FILLCELL_X8 FILLER_82_1202 ();
 FILLCELL_X1 FILLER_82_1216 ();
 FILLCELL_X2 FILLER_82_1236 ();
 FILLCELL_X16 FILLER_83_1 ();
 FILLCELL_X2 FILLER_83_17 ();
 FILLCELL_X1 FILLER_83_24 ();
 FILLCELL_X1 FILLER_83_52 ();
 FILLCELL_X8 FILLER_83_74 ();
 FILLCELL_X4 FILLER_83_82 ();
 FILLCELL_X2 FILLER_83_86 ();
 FILLCELL_X4 FILLER_83_95 ();
 FILLCELL_X2 FILLER_83_126 ();
 FILLCELL_X8 FILLER_83_135 ();
 FILLCELL_X1 FILLER_83_143 ();
 FILLCELL_X16 FILLER_83_164 ();
 FILLCELL_X1 FILLER_83_183 ();
 FILLCELL_X4 FILLER_83_197 ();
 FILLCELL_X2 FILLER_83_201 ();
 FILLCELL_X1 FILLER_83_203 ();
 FILLCELL_X4 FILLER_83_252 ();
 FILLCELL_X2 FILLER_83_256 ();
 FILLCELL_X1 FILLER_83_258 ();
 FILLCELL_X4 FILLER_83_299 ();
 FILLCELL_X1 FILLER_83_303 ();
 FILLCELL_X1 FILLER_83_324 ();
 FILLCELL_X1 FILLER_83_345 ();
 FILLCELL_X1 FILLER_83_349 ();
 FILLCELL_X1 FILLER_83_353 ();
 FILLCELL_X1 FILLER_83_374 ();
 FILLCELL_X2 FILLER_83_392 ();
 FILLCELL_X8 FILLER_83_401 ();
 FILLCELL_X2 FILLER_83_416 ();
 FILLCELL_X4 FILLER_83_438 ();
 FILLCELL_X2 FILLER_83_442 ();
 FILLCELL_X1 FILLER_83_444 ();
 FILLCELL_X1 FILLER_83_454 ();
 FILLCELL_X4 FILLER_83_458 ();
 FILLCELL_X2 FILLER_83_462 ();
 FILLCELL_X8 FILLER_83_471 ();
 FILLCELL_X16 FILLER_83_486 ();
 FILLCELL_X4 FILLER_83_511 ();
 FILLCELL_X4 FILLER_83_528 ();
 FILLCELL_X2 FILLER_83_536 ();
 FILLCELL_X2 FILLER_83_542 ();
 FILLCELL_X8 FILLER_83_579 ();
 FILLCELL_X4 FILLER_83_587 ();
 FILLCELL_X2 FILLER_83_591 ();
 FILLCELL_X1 FILLER_83_593 ();
 FILLCELL_X8 FILLER_83_608 ();
 FILLCELL_X1 FILLER_83_630 ();
 FILLCELL_X2 FILLER_83_640 ();
 FILLCELL_X1 FILLER_83_642 ();
 FILLCELL_X8 FILLER_83_648 ();
 FILLCELL_X4 FILLER_83_656 ();
 FILLCELL_X16 FILLER_83_667 ();
 FILLCELL_X4 FILLER_83_683 ();
 FILLCELL_X2 FILLER_83_687 ();
 FILLCELL_X4 FILLER_83_709 ();
 FILLCELL_X4 FILLER_83_716 ();
 FILLCELL_X16 FILLER_83_724 ();
 FILLCELL_X1 FILLER_83_744 ();
 FILLCELL_X8 FILLER_83_752 ();
 FILLCELL_X1 FILLER_83_760 ();
 FILLCELL_X8 FILLER_83_766 ();
 FILLCELL_X4 FILLER_83_774 ();
 FILLCELL_X2 FILLER_83_782 ();
 FILLCELL_X4 FILLER_83_802 ();
 FILLCELL_X2 FILLER_83_806 ();
 FILLCELL_X16 FILLER_83_813 ();
 FILLCELL_X8 FILLER_83_829 ();
 FILLCELL_X4 FILLER_83_837 ();
 FILLCELL_X1 FILLER_83_841 ();
 FILLCELL_X8 FILLER_83_846 ();
 FILLCELL_X4 FILLER_83_854 ();
 FILLCELL_X8 FILLER_83_868 ();
 FILLCELL_X4 FILLER_83_883 ();
 FILLCELL_X2 FILLER_83_887 ();
 FILLCELL_X1 FILLER_83_889 ();
 FILLCELL_X8 FILLER_83_895 ();
 FILLCELL_X2 FILLER_83_903 ();
 FILLCELL_X1 FILLER_83_933 ();
 FILLCELL_X2 FILLER_83_937 ();
 FILLCELL_X1 FILLER_83_939 ();
 FILLCELL_X2 FILLER_83_947 ();
 FILLCELL_X1 FILLER_83_963 ();
 FILLCELL_X1 FILLER_83_971 ();
 FILLCELL_X4 FILLER_83_983 ();
 FILLCELL_X4 FILLER_83_1002 ();
 FILLCELL_X1 FILLER_83_1037 ();
 FILLCELL_X16 FILLER_83_1045 ();
 FILLCELL_X8 FILLER_83_1061 ();
 FILLCELL_X2 FILLER_83_1069 ();
 FILLCELL_X1 FILLER_83_1071 ();
 FILLCELL_X4 FILLER_83_1079 ();
 FILLCELL_X1 FILLER_83_1083 ();
 FILLCELL_X1 FILLER_83_1087 ();
 FILLCELL_X2 FILLER_83_1095 ();
 FILLCELL_X4 FILLER_83_1104 ();
 FILLCELL_X2 FILLER_83_1134 ();
 FILLCELL_X4 FILLER_83_1141 ();
 FILLCELL_X2 FILLER_83_1145 ();
 FILLCELL_X1 FILLER_83_1147 ();
 FILLCELL_X4 FILLER_83_1153 ();
 FILLCELL_X1 FILLER_83_1157 ();
 FILLCELL_X1 FILLER_83_1166 ();
 FILLCELL_X8 FILLER_83_1171 ();
 FILLCELL_X1 FILLER_83_1179 ();
 FILLCELL_X4 FILLER_83_1208 ();
 FILLCELL_X1 FILLER_83_1212 ();
 FILLCELL_X4 FILLER_83_1217 ();
 FILLCELL_X1 FILLER_83_1221 ();
 FILLCELL_X2 FILLER_83_1235 ();
 FILLCELL_X2 FILLER_83_1250 ();
 FILLCELL_X1 FILLER_84_1 ();
 FILLCELL_X4 FILLER_84_22 ();
 FILLCELL_X2 FILLER_84_26 ();
 FILLCELL_X1 FILLER_84_28 ();
 FILLCELL_X4 FILLER_84_36 ();
 FILLCELL_X2 FILLER_84_40 ();
 FILLCELL_X1 FILLER_84_42 ();
 FILLCELL_X8 FILLER_84_70 ();
 FILLCELL_X4 FILLER_84_78 ();
 FILLCELL_X8 FILLER_84_102 ();
 FILLCELL_X2 FILLER_84_110 ();
 FILLCELL_X8 FILLER_84_119 ();
 FILLCELL_X1 FILLER_84_157 ();
 FILLCELL_X1 FILLER_84_165 ();
 FILLCELL_X8 FILLER_84_192 ();
 FILLCELL_X8 FILLER_84_207 ();
 FILLCELL_X4 FILLER_84_227 ();
 FILLCELL_X2 FILLER_84_231 ();
 FILLCELL_X1 FILLER_84_233 ();
 FILLCELL_X2 FILLER_84_255 ();
 FILLCELL_X1 FILLER_84_257 ();
 FILLCELL_X2 FILLER_84_288 ();
 FILLCELL_X8 FILLER_84_307 ();
 FILLCELL_X8 FILLER_84_317 ();
 FILLCELL_X2 FILLER_84_325 ();
 FILLCELL_X1 FILLER_84_327 ();
 FILLCELL_X4 FILLER_84_331 ();
 FILLCELL_X2 FILLER_84_335 ();
 FILLCELL_X2 FILLER_84_344 ();
 FILLCELL_X4 FILLER_84_393 ();
 FILLCELL_X2 FILLER_84_397 ();
 FILLCELL_X16 FILLER_84_410 ();
 FILLCELL_X1 FILLER_84_426 ();
 FILLCELL_X2 FILLER_84_434 ();
 FILLCELL_X4 FILLER_84_446 ();
 FILLCELL_X2 FILLER_84_450 ();
 FILLCELL_X1 FILLER_84_452 ();
 FILLCELL_X4 FILLER_84_457 ();
 FILLCELL_X8 FILLER_84_464 ();
 FILLCELL_X8 FILLER_84_479 ();
 FILLCELL_X4 FILLER_84_487 ();
 FILLCELL_X4 FILLER_84_518 ();
 FILLCELL_X2 FILLER_84_522 ();
 FILLCELL_X1 FILLER_84_524 ();
 FILLCELL_X1 FILLER_84_560 ();
 FILLCELL_X8 FILLER_84_568 ();
 FILLCELL_X4 FILLER_84_576 ();
 FILLCELL_X2 FILLER_84_580 ();
 FILLCELL_X1 FILLER_84_582 ();
 FILLCELL_X4 FILLER_84_616 ();
 FILLCELL_X8 FILLER_84_623 ();
 FILLCELL_X8 FILLER_84_632 ();
 FILLCELL_X4 FILLER_84_640 ();
 FILLCELL_X1 FILLER_84_644 ();
 FILLCELL_X2 FILLER_84_661 ();
 FILLCELL_X1 FILLER_84_663 ();
 FILLCELL_X1 FILLER_84_691 ();
 FILLCELL_X1 FILLER_84_702 ();
 FILLCELL_X1 FILLER_84_707 ();
 FILLCELL_X1 FILLER_84_722 ();
 FILLCELL_X8 FILLER_84_730 ();
 FILLCELL_X1 FILLER_84_754 ();
 FILLCELL_X8 FILLER_84_760 ();
 FILLCELL_X1 FILLER_84_768 ();
 FILLCELL_X1 FILLER_84_779 ();
 FILLCELL_X8 FILLER_84_789 ();
 FILLCELL_X1 FILLER_84_797 ();
 FILLCELL_X4 FILLER_84_804 ();
 FILLCELL_X1 FILLER_84_808 ();
 FILLCELL_X4 FILLER_84_836 ();
 FILLCELL_X1 FILLER_84_840 ();
 FILLCELL_X4 FILLER_84_851 ();
 FILLCELL_X4 FILLER_84_873 ();
 FILLCELL_X16 FILLER_84_901 ();
 FILLCELL_X4 FILLER_84_917 ();
 FILLCELL_X2 FILLER_84_921 ();
 FILLCELL_X1 FILLER_84_934 ();
 FILLCELL_X2 FILLER_84_938 ();
 FILLCELL_X4 FILLER_84_960 ();
 FILLCELL_X8 FILLER_84_966 ();
 FILLCELL_X2 FILLER_84_974 ();
 FILLCELL_X8 FILLER_84_985 ();
 FILLCELL_X1 FILLER_84_993 ();
 FILLCELL_X2 FILLER_84_997 ();
 FILLCELL_X2 FILLER_84_1021 ();
 FILLCELL_X1 FILLER_84_1023 ();
 FILLCELL_X2 FILLER_84_1030 ();
 FILLCELL_X2 FILLER_84_1035 ();
 FILLCELL_X4 FILLER_84_1053 ();
 FILLCELL_X2 FILLER_84_1085 ();
 FILLCELL_X2 FILLER_84_1112 ();
 FILLCELL_X2 FILLER_84_1126 ();
 FILLCELL_X1 FILLER_84_1128 ();
 FILLCELL_X4 FILLER_84_1138 ();
 FILLCELL_X1 FILLER_84_1142 ();
 FILLCELL_X4 FILLER_84_1177 ();
 FILLCELL_X2 FILLER_84_1181 ();
 FILLCELL_X2 FILLER_84_1206 ();
 FILLCELL_X2 FILLER_84_1228 ();
 FILLCELL_X8 FILLER_85_1 ();
 FILLCELL_X4 FILLER_85_9 ();
 FILLCELL_X16 FILLER_85_47 ();
 FILLCELL_X4 FILLER_85_63 ();
 FILLCELL_X2 FILLER_85_67 ();
 FILLCELL_X4 FILLER_85_76 ();
 FILLCELL_X2 FILLER_85_80 ();
 FILLCELL_X1 FILLER_85_101 ();
 FILLCELL_X8 FILLER_85_109 ();
 FILLCELL_X2 FILLER_85_117 ();
 FILLCELL_X1 FILLER_85_126 ();
 FILLCELL_X4 FILLER_85_134 ();
 FILLCELL_X2 FILLER_85_138 ();
 FILLCELL_X1 FILLER_85_147 ();
 FILLCELL_X2 FILLER_85_156 ();
 FILLCELL_X1 FILLER_85_158 ();
 FILLCELL_X4 FILLER_85_179 ();
 FILLCELL_X1 FILLER_85_183 ();
 FILLCELL_X4 FILLER_85_191 ();
 FILLCELL_X2 FILLER_85_195 ();
 FILLCELL_X1 FILLER_85_197 ();
 FILLCELL_X4 FILLER_85_205 ();
 FILLCELL_X1 FILLER_85_229 ();
 FILLCELL_X4 FILLER_85_237 ();
 FILLCELL_X1 FILLER_85_241 ();
 FILLCELL_X8 FILLER_85_249 ();
 FILLCELL_X4 FILLER_85_257 ();
 FILLCELL_X4 FILLER_85_269 ();
 FILLCELL_X8 FILLER_85_276 ();
 FILLCELL_X1 FILLER_85_295 ();
 FILLCELL_X4 FILLER_85_299 ();
 FILLCELL_X2 FILLER_85_303 ();
 FILLCELL_X1 FILLER_85_309 ();
 FILLCELL_X8 FILLER_85_332 ();
 FILLCELL_X32 FILLER_85_360 ();
 FILLCELL_X1 FILLER_85_405 ();
 FILLCELL_X4 FILLER_85_433 ();
 FILLCELL_X1 FILLER_85_437 ();
 FILLCELL_X4 FILLER_85_470 ();
 FILLCELL_X2 FILLER_85_481 ();
 FILLCELL_X2 FILLER_85_503 ();
 FILLCELL_X4 FILLER_85_508 ();
 FILLCELL_X1 FILLER_85_512 ();
 FILLCELL_X2 FILLER_85_532 ();
 FILLCELL_X1 FILLER_85_534 ();
 FILLCELL_X16 FILLER_85_572 ();
 FILLCELL_X2 FILLER_85_588 ();
 FILLCELL_X1 FILLER_85_590 ();
 FILLCELL_X1 FILLER_85_595 ();
 FILLCELL_X2 FILLER_85_599 ();
 FILLCELL_X8 FILLER_85_608 ();
 FILLCELL_X2 FILLER_85_616 ();
 FILLCELL_X1 FILLER_85_618 ();
 FILLCELL_X2 FILLER_85_637 ();
 FILLCELL_X1 FILLER_85_639 ();
 FILLCELL_X4 FILLER_85_654 ();
 FILLCELL_X1 FILLER_85_658 ();
 FILLCELL_X4 FILLER_85_677 ();
 FILLCELL_X2 FILLER_85_681 ();
 FILLCELL_X1 FILLER_85_683 ();
 FILLCELL_X1 FILLER_85_709 ();
 FILLCELL_X1 FILLER_85_726 ();
 FILLCELL_X4 FILLER_85_746 ();
 FILLCELL_X1 FILLER_85_759 ();
 FILLCELL_X8 FILLER_85_763 ();
 FILLCELL_X4 FILLER_85_771 ();
 FILLCELL_X2 FILLER_85_794 ();
 FILLCELL_X1 FILLER_85_796 ();
 FILLCELL_X8 FILLER_85_808 ();
 FILLCELL_X2 FILLER_85_816 ();
 FILLCELL_X1 FILLER_85_818 ();
 FILLCELL_X8 FILLER_85_822 ();
 FILLCELL_X4 FILLER_85_830 ();
 FILLCELL_X1 FILLER_85_834 ();
 FILLCELL_X4 FILLER_85_839 ();
 FILLCELL_X2 FILLER_85_843 ();
 FILLCELL_X1 FILLER_85_845 ();
 FILLCELL_X16 FILLER_85_854 ();
 FILLCELL_X4 FILLER_85_870 ();
 FILLCELL_X8 FILLER_85_898 ();
 FILLCELL_X1 FILLER_85_906 ();
 FILLCELL_X1 FILLER_85_921 ();
 FILLCELL_X2 FILLER_85_926 ();
 FILLCELL_X1 FILLER_85_952 ();
 FILLCELL_X2 FILLER_85_960 ();
 FILLCELL_X2 FILLER_85_969 ();
 FILLCELL_X8 FILLER_85_985 ();
 FILLCELL_X16 FILLER_85_1001 ();
 FILLCELL_X2 FILLER_85_1017 ();
 FILLCELL_X1 FILLER_85_1019 ();
 FILLCELL_X4 FILLER_85_1024 ();
 FILLCELL_X1 FILLER_85_1028 ();
 FILLCELL_X1 FILLER_85_1059 ();
 FILLCELL_X1 FILLER_85_1067 ();
 FILLCELL_X1 FILLER_85_1081 ();
 FILLCELL_X1 FILLER_85_1089 ();
 FILLCELL_X2 FILLER_85_1107 ();
 FILLCELL_X2 FILLER_85_1130 ();
 FILLCELL_X8 FILLER_85_1139 ();
 FILLCELL_X1 FILLER_85_1161 ();
 FILLCELL_X4 FILLER_85_1167 ();
 FILLCELL_X2 FILLER_85_1171 ();
 FILLCELL_X1 FILLER_85_1173 ();
 FILLCELL_X4 FILLER_85_1178 ();
 FILLCELL_X1 FILLER_85_1196 ();
 FILLCELL_X2 FILLER_85_1211 ();
 FILLCELL_X4 FILLER_85_1218 ();
 FILLCELL_X2 FILLER_85_1222 ();
 FILLCELL_X4 FILLER_85_1251 ();
 FILLCELL_X16 FILLER_86_1 ();
 FILLCELL_X4 FILLER_86_17 ();
 FILLCELL_X1 FILLER_86_21 ();
 FILLCELL_X16 FILLER_86_36 ();
 FILLCELL_X2 FILLER_86_52 ();
 FILLCELL_X1 FILLER_86_54 ();
 FILLCELL_X8 FILLER_86_62 ();
 FILLCELL_X4 FILLER_86_70 ();
 FILLCELL_X1 FILLER_86_74 ();
 FILLCELL_X2 FILLER_86_95 ();
 FILLCELL_X1 FILLER_86_97 ();
 FILLCELL_X16 FILLER_86_139 ();
 FILLCELL_X4 FILLER_86_155 ();
 FILLCELL_X8 FILLER_86_179 ();
 FILLCELL_X4 FILLER_86_187 ();
 FILLCELL_X1 FILLER_86_204 ();
 FILLCELL_X1 FILLER_86_228 ();
 FILLCELL_X1 FILLER_86_236 ();
 FILLCELL_X1 FILLER_86_251 ();
 FILLCELL_X2 FILLER_86_255 ();
 FILLCELL_X2 FILLER_86_271 ();
 FILLCELL_X1 FILLER_86_307 ();
 FILLCELL_X2 FILLER_86_321 ();
 FILLCELL_X16 FILLER_86_344 ();
 FILLCELL_X1 FILLER_86_360 ();
 FILLCELL_X1 FILLER_86_366 ();
 FILLCELL_X4 FILLER_86_377 ();
 FILLCELL_X2 FILLER_86_385 ();
 FILLCELL_X8 FILLER_86_390 ();
 FILLCELL_X2 FILLER_86_398 ();
 FILLCELL_X1 FILLER_86_400 ();
 FILLCELL_X2 FILLER_86_405 ();
 FILLCELL_X1 FILLER_86_407 ();
 FILLCELL_X4 FILLER_86_432 ();
 FILLCELL_X2 FILLER_86_436 ();
 FILLCELL_X2 FILLER_86_442 ();
 FILLCELL_X2 FILLER_86_447 ();
 FILLCELL_X4 FILLER_86_469 ();
 FILLCELL_X1 FILLER_86_493 ();
 FILLCELL_X1 FILLER_86_501 ();
 FILLCELL_X2 FILLER_86_509 ();
 FILLCELL_X8 FILLER_86_521 ();
 FILLCELL_X4 FILLER_86_529 ();
 FILLCELL_X8 FILLER_86_563 ();
 FILLCELL_X4 FILLER_86_578 ();
 FILLCELL_X1 FILLER_86_609 ();
 FILLCELL_X8 FILLER_86_617 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X8 FILLER_86_632 ();
 FILLCELL_X4 FILLER_86_640 ();
 FILLCELL_X2 FILLER_86_644 ();
 FILLCELL_X8 FILLER_86_660 ();
 FILLCELL_X2 FILLER_86_673 ();
 FILLCELL_X8 FILLER_86_678 ();
 FILLCELL_X4 FILLER_86_686 ();
 FILLCELL_X2 FILLER_86_690 ();
 FILLCELL_X1 FILLER_86_692 ();
 FILLCELL_X4 FILLER_86_702 ();
 FILLCELL_X2 FILLER_86_706 ();
 FILLCELL_X1 FILLER_86_708 ();
 FILLCELL_X8 FILLER_86_713 ();
 FILLCELL_X1 FILLER_86_721 ();
 FILLCELL_X4 FILLER_86_732 ();
 FILLCELL_X4 FILLER_86_766 ();
 FILLCELL_X2 FILLER_86_773 ();
 FILLCELL_X1 FILLER_86_775 ();
 FILLCELL_X4 FILLER_86_785 ();
 FILLCELL_X2 FILLER_86_789 ();
 FILLCELL_X8 FILLER_86_798 ();
 FILLCELL_X2 FILLER_86_806 ();
 FILLCELL_X8 FILLER_86_819 ();
 FILLCELL_X2 FILLER_86_827 ();
 FILLCELL_X8 FILLER_86_857 ();
 FILLCELL_X1 FILLER_86_868 ();
 FILLCELL_X1 FILLER_86_883 ();
 FILLCELL_X8 FILLER_86_892 ();
 FILLCELL_X4 FILLER_86_900 ();
 FILLCELL_X4 FILLER_86_913 ();
 FILLCELL_X2 FILLER_86_917 ();
 FILLCELL_X1 FILLER_86_949 ();
 FILLCELL_X1 FILLER_86_964 ();
 FILLCELL_X1 FILLER_86_989 ();
 FILLCELL_X4 FILLER_86_1005 ();
 FILLCELL_X2 FILLER_86_1009 ();
 FILLCELL_X1 FILLER_86_1011 ();
 FILLCELL_X2 FILLER_86_1031 ();
 FILLCELL_X1 FILLER_86_1033 ();
 FILLCELL_X2 FILLER_86_1041 ();
 FILLCELL_X4 FILLER_86_1050 ();
 FILLCELL_X2 FILLER_86_1061 ();
 FILLCELL_X1 FILLER_86_1063 ();
 FILLCELL_X8 FILLER_86_1074 ();
 FILLCELL_X2 FILLER_86_1082 ();
 FILLCELL_X16 FILLER_86_1115 ();
 FILLCELL_X8 FILLER_86_1161 ();
 FILLCELL_X4 FILLER_86_1169 ();
 FILLCELL_X1 FILLER_86_1179 ();
 FILLCELL_X2 FILLER_86_1184 ();
 FILLCELL_X2 FILLER_86_1190 ();
 FILLCELL_X1 FILLER_86_1192 ();
 FILLCELL_X8 FILLER_86_1199 ();
 FILLCELL_X4 FILLER_86_1207 ();
 FILLCELL_X1 FILLER_86_1211 ();
 FILLCELL_X4 FILLER_86_1216 ();
 FILLCELL_X2 FILLER_86_1220 ();
 FILLCELL_X1 FILLER_86_1229 ();
 FILLCELL_X2 FILLER_86_1233 ();
 FILLCELL_X4 FILLER_86_1238 ();
 FILLCELL_X4 FILLER_86_1249 ();
 FILLCELL_X2 FILLER_86_1253 ();
 FILLCELL_X2 FILLER_87_1 ();
 FILLCELL_X4 FILLER_87_23 ();
 FILLCELL_X1 FILLER_87_27 ();
 FILLCELL_X8 FILLER_87_35 ();
 FILLCELL_X2 FILLER_87_43 ();
 FILLCELL_X2 FILLER_87_65 ();
 FILLCELL_X1 FILLER_87_67 ();
 FILLCELL_X4 FILLER_87_116 ();
 FILLCELL_X2 FILLER_87_120 ();
 FILLCELL_X4 FILLER_87_170 ();
 FILLCELL_X2 FILLER_87_174 ();
 FILLCELL_X1 FILLER_87_176 ();
 FILLCELL_X1 FILLER_87_192 ();
 FILLCELL_X8 FILLER_87_200 ();
 FILLCELL_X2 FILLER_87_208 ();
 FILLCELL_X8 FILLER_87_224 ();
 FILLCELL_X1 FILLER_87_232 ();
 FILLCELL_X8 FILLER_87_247 ();
 FILLCELL_X4 FILLER_87_255 ();
 FILLCELL_X4 FILLER_87_282 ();
 FILLCELL_X1 FILLER_87_286 ();
 FILLCELL_X1 FILLER_87_294 ();
 FILLCELL_X1 FILLER_87_302 ();
 FILLCELL_X1 FILLER_87_306 ();
 FILLCELL_X4 FILLER_87_310 ();
 FILLCELL_X4 FILLER_87_318 ();
 FILLCELL_X1 FILLER_87_322 ();
 FILLCELL_X8 FILLER_87_326 ();
 FILLCELL_X4 FILLER_87_334 ();
 FILLCELL_X1 FILLER_87_352 ();
 FILLCELL_X8 FILLER_87_413 ();
 FILLCELL_X4 FILLER_87_426 ();
 FILLCELL_X2 FILLER_87_430 ();
 FILLCELL_X1 FILLER_87_432 ();
 FILLCELL_X1 FILLER_87_453 ();
 FILLCELL_X2 FILLER_87_461 ();
 FILLCELL_X1 FILLER_87_463 ();
 FILLCELL_X16 FILLER_87_478 ();
 FILLCELL_X4 FILLER_87_494 ();
 FILLCELL_X2 FILLER_87_498 ();
 FILLCELL_X8 FILLER_87_539 ();
 FILLCELL_X1 FILLER_87_547 ();
 FILLCELL_X8 FILLER_87_572 ();
 FILLCELL_X2 FILLER_87_580 ();
 FILLCELL_X1 FILLER_87_582 ();
 FILLCELL_X4 FILLER_87_590 ();
 FILLCELL_X4 FILLER_87_615 ();
 FILLCELL_X16 FILLER_87_637 ();
 FILLCELL_X2 FILLER_87_653 ();
 FILLCELL_X8 FILLER_87_662 ();
 FILLCELL_X4 FILLER_87_670 ();
 FILLCELL_X1 FILLER_87_674 ();
 FILLCELL_X16 FILLER_87_684 ();
 FILLCELL_X8 FILLER_87_700 ();
 FILLCELL_X8 FILLER_87_721 ();
 FILLCELL_X2 FILLER_87_729 ();
 FILLCELL_X2 FILLER_87_745 ();
 FILLCELL_X1 FILLER_87_747 ();
 FILLCELL_X2 FILLER_87_768 ();
 FILLCELL_X1 FILLER_87_784 ();
 FILLCELL_X1 FILLER_87_795 ();
 FILLCELL_X2 FILLER_87_807 ();
 FILLCELL_X1 FILLER_87_809 ();
 FILLCELL_X8 FILLER_87_817 ();
 FILLCELL_X2 FILLER_87_825 ();
 FILLCELL_X4 FILLER_87_834 ();
 FILLCELL_X2 FILLER_87_838 ();
 FILLCELL_X2 FILLER_87_869 ();
 FILLCELL_X1 FILLER_87_871 ();
 FILLCELL_X1 FILLER_87_891 ();
 FILLCELL_X8 FILLER_87_902 ();
 FILLCELL_X2 FILLER_87_910 ();
 FILLCELL_X1 FILLER_87_912 ();
 FILLCELL_X4 FILLER_87_923 ();
 FILLCELL_X1 FILLER_87_927 ();
 FILLCELL_X1 FILLER_87_939 ();
 FILLCELL_X1 FILLER_87_951 ();
 FILLCELL_X2 FILLER_87_1013 ();
 FILLCELL_X8 FILLER_87_1019 ();
 FILLCELL_X4 FILLER_87_1027 ();
 FILLCELL_X1 FILLER_87_1031 ();
 FILLCELL_X1 FILLER_87_1043 ();
 FILLCELL_X8 FILLER_87_1058 ();
 FILLCELL_X2 FILLER_87_1072 ();
 FILLCELL_X1 FILLER_87_1074 ();
 FILLCELL_X2 FILLER_87_1082 ();
 FILLCELL_X1 FILLER_87_1084 ();
 FILLCELL_X16 FILLER_87_1092 ();
 FILLCELL_X2 FILLER_87_1108 ();
 FILLCELL_X1 FILLER_87_1110 ();
 FILLCELL_X16 FILLER_87_1116 ();
 FILLCELL_X2 FILLER_87_1132 ();
 FILLCELL_X4 FILLER_87_1145 ();
 FILLCELL_X2 FILLER_87_1149 ();
 FILLCELL_X8 FILLER_87_1156 ();
 FILLCELL_X4 FILLER_87_1164 ();
 FILLCELL_X2 FILLER_87_1198 ();
 FILLCELL_X4 FILLER_87_1217 ();
 FILLCELL_X2 FILLER_87_1221 ();
 FILLCELL_X1 FILLER_87_1223 ();
 FILLCELL_X1 FILLER_87_1230 ();
 FILLCELL_X8 FILLER_88_1 ();
 FILLCELL_X2 FILLER_88_9 ();
 FILLCELL_X1 FILLER_88_11 ();
 FILLCELL_X4 FILLER_88_19 ();
 FILLCELL_X2 FILLER_88_23 ();
 FILLCELL_X1 FILLER_88_32 ();
 FILLCELL_X1 FILLER_88_47 ();
 FILLCELL_X2 FILLER_88_55 ();
 FILLCELL_X2 FILLER_88_84 ();
 FILLCELL_X1 FILLER_88_86 ();
 FILLCELL_X2 FILLER_88_94 ();
 FILLCELL_X1 FILLER_88_96 ();
 FILLCELL_X2 FILLER_88_111 ();
 FILLCELL_X1 FILLER_88_140 ();
 FILLCELL_X8 FILLER_88_148 ();
 FILLCELL_X2 FILLER_88_176 ();
 FILLCELL_X8 FILLER_88_181 ();
 FILLCELL_X2 FILLER_88_202 ();
 FILLCELL_X1 FILLER_88_204 ();
 FILLCELL_X1 FILLER_88_225 ();
 FILLCELL_X16 FILLER_88_240 ();
 FILLCELL_X2 FILLER_88_256 ();
 FILLCELL_X1 FILLER_88_258 ();
 FILLCELL_X2 FILLER_88_270 ();
 FILLCELL_X4 FILLER_88_332 ();
 FILLCELL_X1 FILLER_88_336 ();
 FILLCELL_X4 FILLER_88_351 ();
 FILLCELL_X2 FILLER_88_355 ();
 FILLCELL_X1 FILLER_88_357 ();
 FILLCELL_X1 FILLER_88_364 ();
 FILLCELL_X4 FILLER_88_377 ();
 FILLCELL_X2 FILLER_88_381 ();
 FILLCELL_X2 FILLER_88_387 ();
 FILLCELL_X8 FILLER_88_392 ();
 FILLCELL_X2 FILLER_88_400 ();
 FILLCELL_X8 FILLER_88_433 ();
 FILLCELL_X2 FILLER_88_441 ();
 FILLCELL_X1 FILLER_88_443 ();
 FILLCELL_X16 FILLER_88_516 ();
 FILLCELL_X4 FILLER_88_566 ();
 FILLCELL_X1 FILLER_88_570 ();
 FILLCELL_X2 FILLER_88_585 ();
 FILLCELL_X1 FILLER_88_587 ();
 FILLCELL_X2 FILLER_88_628 ();
 FILLCELL_X1 FILLER_88_630 ();
 FILLCELL_X2 FILLER_88_636 ();
 FILLCELL_X1 FILLER_88_638 ();
 FILLCELL_X16 FILLER_88_642 ();
 FILLCELL_X4 FILLER_88_658 ();
 FILLCELL_X2 FILLER_88_662 ();
 FILLCELL_X1 FILLER_88_664 ();
 FILLCELL_X1 FILLER_88_679 ();
 FILLCELL_X8 FILLER_88_701 ();
 FILLCELL_X4 FILLER_88_709 ();
 FILLCELL_X1 FILLER_88_713 ();
 FILLCELL_X8 FILLER_88_721 ();
 FILLCELL_X4 FILLER_88_729 ();
 FILLCELL_X2 FILLER_88_733 ();
 FILLCELL_X16 FILLER_88_742 ();
 FILLCELL_X2 FILLER_88_758 ();
 FILLCELL_X4 FILLER_88_771 ();
 FILLCELL_X1 FILLER_88_775 ();
 FILLCELL_X4 FILLER_88_781 ();
 FILLCELL_X2 FILLER_88_785 ();
 FILLCELL_X1 FILLER_88_794 ();
 FILLCELL_X16 FILLER_88_803 ();
 FILLCELL_X8 FILLER_88_819 ();
 FILLCELL_X2 FILLER_88_827 ();
 FILLCELL_X1 FILLER_88_846 ();
 FILLCELL_X2 FILLER_88_858 ();
 FILLCELL_X4 FILLER_88_882 ();
 FILLCELL_X2 FILLER_88_903 ();
 FILLCELL_X2 FILLER_88_909 ();
 FILLCELL_X4 FILLER_88_932 ();
 FILLCELL_X1 FILLER_88_936 ();
 FILLCELL_X8 FILLER_88_951 ();
 FILLCELL_X8 FILLER_88_966 ();
 FILLCELL_X4 FILLER_88_974 ();
 FILLCELL_X2 FILLER_88_978 ();
 FILLCELL_X1 FILLER_88_980 ();
 FILLCELL_X2 FILLER_88_995 ();
 FILLCELL_X1 FILLER_88_997 ();
 FILLCELL_X8 FILLER_88_1001 ();
 FILLCELL_X4 FILLER_88_1009 ();
 FILLCELL_X2 FILLER_88_1013 ();
 FILLCELL_X1 FILLER_88_1046 ();
 FILLCELL_X1 FILLER_88_1084 ();
 FILLCELL_X8 FILLER_88_1092 ();
 FILLCELL_X1 FILLER_88_1100 ();
 FILLCELL_X8 FILLER_88_1128 ();
 FILLCELL_X4 FILLER_88_1162 ();
 FILLCELL_X2 FILLER_88_1166 ();
 FILLCELL_X8 FILLER_88_1209 ();
 FILLCELL_X4 FILLER_88_1217 ();
 FILLCELL_X1 FILLER_88_1221 ();
 FILLCELL_X4 FILLER_88_1229 ();
 FILLCELL_X2 FILLER_88_1233 ();
 FILLCELL_X1 FILLER_88_1235 ();
 FILLCELL_X8 FILLER_88_1243 ();
 FILLCELL_X4 FILLER_88_1251 ();
 FILLCELL_X1 FILLER_89_1 ();
 FILLCELL_X2 FILLER_89_29 ();
 FILLCELL_X8 FILLER_89_46 ();
 FILLCELL_X4 FILLER_89_81 ();
 FILLCELL_X2 FILLER_89_92 ();
 FILLCELL_X1 FILLER_89_94 ();
 FILLCELL_X4 FILLER_89_102 ();
 FILLCELL_X2 FILLER_89_106 ();
 FILLCELL_X1 FILLER_89_108 ();
 FILLCELL_X2 FILLER_89_123 ();
 FILLCELL_X8 FILLER_89_139 ();
 FILLCELL_X4 FILLER_89_147 ();
 FILLCELL_X2 FILLER_89_151 ();
 FILLCELL_X2 FILLER_89_156 ();
 FILLCELL_X1 FILLER_89_165 ();
 FILLCELL_X2 FILLER_89_171 ();
 FILLCELL_X8 FILLER_89_179 ();
 FILLCELL_X4 FILLER_89_187 ();
 FILLCELL_X2 FILLER_89_194 ();
 FILLCELL_X1 FILLER_89_196 ();
 FILLCELL_X2 FILLER_89_204 ();
 FILLCELL_X1 FILLER_89_206 ();
 FILLCELL_X2 FILLER_89_218 ();
 FILLCELL_X1 FILLER_89_220 ();
 FILLCELL_X4 FILLER_89_241 ();
 FILLCELL_X1 FILLER_89_245 ();
 FILLCELL_X4 FILLER_89_253 ();
 FILLCELL_X2 FILLER_89_257 ();
 FILLCELL_X1 FILLER_89_259 ();
 FILLCELL_X16 FILLER_89_283 ();
 FILLCELL_X4 FILLER_89_299 ();
 FILLCELL_X2 FILLER_89_303 ();
 FILLCELL_X16 FILLER_89_311 ();
 FILLCELL_X4 FILLER_89_327 ();
 FILLCELL_X2 FILLER_89_331 ();
 FILLCELL_X2 FILLER_89_353 ();
 FILLCELL_X4 FILLER_89_375 ();
 FILLCELL_X1 FILLER_89_403 ();
 FILLCELL_X8 FILLER_89_407 ();
 FILLCELL_X8 FILLER_89_422 ();
 FILLCELL_X2 FILLER_89_430 ();
 FILLCELL_X1 FILLER_89_432 ();
 FILLCELL_X8 FILLER_89_453 ();
 FILLCELL_X4 FILLER_89_477 ();
 FILLCELL_X2 FILLER_89_481 ();
 FILLCELL_X8 FILLER_89_492 ();
 FILLCELL_X4 FILLER_89_500 ();
 FILLCELL_X2 FILLER_89_504 ();
 FILLCELL_X8 FILLER_89_523 ();
 FILLCELL_X2 FILLER_89_531 ();
 FILLCELL_X4 FILLER_89_582 ();
 FILLCELL_X1 FILLER_89_586 ();
 FILLCELL_X1 FILLER_89_609 ();
 FILLCELL_X8 FILLER_89_617 ();
 FILLCELL_X4 FILLER_89_625 ();
 FILLCELL_X2 FILLER_89_629 ();
 FILLCELL_X1 FILLER_89_631 ();
 FILLCELL_X4 FILLER_89_636 ();
 FILLCELL_X1 FILLER_89_645 ();
 FILLCELL_X2 FILLER_89_656 ();
 FILLCELL_X2 FILLER_89_663 ();
 FILLCELL_X1 FILLER_89_672 ();
 FILLCELL_X8 FILLER_89_701 ();
 FILLCELL_X4 FILLER_89_724 ();
 FILLCELL_X2 FILLER_89_728 ();
 FILLCELL_X1 FILLER_89_730 ();
 FILLCELL_X4 FILLER_89_736 ();
 FILLCELL_X2 FILLER_89_740 ();
 FILLCELL_X1 FILLER_89_742 ();
 FILLCELL_X4 FILLER_89_750 ();
 FILLCELL_X1 FILLER_89_754 ();
 FILLCELL_X2 FILLER_89_760 ();
 FILLCELL_X1 FILLER_89_762 ();
 FILLCELL_X4 FILLER_89_767 ();
 FILLCELL_X2 FILLER_89_778 ();
 FILLCELL_X1 FILLER_89_780 ();
 FILLCELL_X2 FILLER_89_784 ();
 FILLCELL_X1 FILLER_89_786 ();
 FILLCELL_X16 FILLER_89_797 ();
 FILLCELL_X4 FILLER_89_820 ();
 FILLCELL_X2 FILLER_89_824 ();
 FILLCELL_X1 FILLER_89_839 ();
 FILLCELL_X2 FILLER_89_846 ();
 FILLCELL_X8 FILLER_89_852 ();
 FILLCELL_X4 FILLER_89_860 ();
 FILLCELL_X1 FILLER_89_867 ();
 FILLCELL_X4 FILLER_89_882 ();
 FILLCELL_X1 FILLER_89_886 ();
 FILLCELL_X1 FILLER_89_904 ();
 FILLCELL_X2 FILLER_89_915 ();
 FILLCELL_X2 FILLER_89_920 ();
 FILLCELL_X4 FILLER_89_942 ();
 FILLCELL_X16 FILLER_89_953 ();
 FILLCELL_X8 FILLER_89_996 ();
 FILLCELL_X1 FILLER_89_1004 ();
 FILLCELL_X8 FILLER_89_1020 ();
 FILLCELL_X4 FILLER_89_1028 ();
 FILLCELL_X2 FILLER_89_1032 ();
 FILLCELL_X1 FILLER_89_1034 ();
 FILLCELL_X1 FILLER_89_1052 ();
 FILLCELL_X4 FILLER_89_1077 ();
 FILLCELL_X4 FILLER_89_1088 ();
 FILLCELL_X2 FILLER_89_1092 ();
 FILLCELL_X2 FILLER_89_1103 ();
 FILLCELL_X1 FILLER_89_1105 ();
 FILLCELL_X1 FILLER_89_1110 ();
 FILLCELL_X2 FILLER_89_1125 ();
 FILLCELL_X1 FILLER_89_1127 ();
 FILLCELL_X2 FILLER_89_1137 ();
 FILLCELL_X4 FILLER_89_1143 ();
 FILLCELL_X2 FILLER_89_1147 ();
 FILLCELL_X8 FILLER_89_1180 ();
 FILLCELL_X4 FILLER_89_1188 ();
 FILLCELL_X2 FILLER_89_1192 ();
 FILLCELL_X1 FILLER_89_1194 ();
 FILLCELL_X1 FILLER_89_1198 ();
 FILLCELL_X8 FILLER_89_1205 ();
 FILLCELL_X2 FILLER_89_1213 ();
 FILLCELL_X4 FILLER_89_1232 ();
 FILLCELL_X4 FILLER_90_1 ();
 FILLCELL_X2 FILLER_90_5 ();
 FILLCELL_X1 FILLER_90_7 ();
 FILLCELL_X8 FILLER_90_42 ();
 FILLCELL_X2 FILLER_90_50 ();
 FILLCELL_X4 FILLER_90_59 ();
 FILLCELL_X2 FILLER_90_63 ();
 FILLCELL_X1 FILLER_90_106 ();
 FILLCELL_X4 FILLER_90_155 ();
 FILLCELL_X2 FILLER_90_159 ();
 FILLCELL_X1 FILLER_90_161 ();
 FILLCELL_X8 FILLER_90_175 ();
 FILLCELL_X1 FILLER_90_183 ();
 FILLCELL_X8 FILLER_90_195 ();
 FILLCELL_X8 FILLER_90_224 ();
 FILLCELL_X4 FILLER_90_232 ();
 FILLCELL_X2 FILLER_90_236 ();
 FILLCELL_X16 FILLER_90_245 ();
 FILLCELL_X2 FILLER_90_261 ();
 FILLCELL_X1 FILLER_90_263 ();
 FILLCELL_X1 FILLER_90_268 ();
 FILLCELL_X1 FILLER_90_273 ();
 FILLCELL_X1 FILLER_90_288 ();
 FILLCELL_X4 FILLER_90_303 ();
 FILLCELL_X16 FILLER_90_331 ();
 FILLCELL_X8 FILLER_90_347 ();
 FILLCELL_X1 FILLER_90_355 ();
 FILLCELL_X4 FILLER_90_365 ();
 FILLCELL_X16 FILLER_90_428 ();
 FILLCELL_X1 FILLER_90_448 ();
 FILLCELL_X4 FILLER_90_452 ();
 FILLCELL_X4 FILLER_90_463 ();
 FILLCELL_X2 FILLER_90_467 ();
 FILLCELL_X4 FILLER_90_487 ();
 FILLCELL_X2 FILLER_90_491 ();
 FILLCELL_X16 FILLER_90_513 ();
 FILLCELL_X1 FILLER_90_529 ();
 FILLCELL_X4 FILLER_90_550 ();
 FILLCELL_X4 FILLER_90_581 ();
 FILLCELL_X2 FILLER_90_585 ();
 FILLCELL_X1 FILLER_90_587 ();
 FILLCELL_X4 FILLER_90_595 ();
 FILLCELL_X2 FILLER_90_599 ();
 FILLCELL_X2 FILLER_90_621 ();
 FILLCELL_X1 FILLER_90_623 ();
 FILLCELL_X2 FILLER_90_641 ();
 FILLCELL_X4 FILLER_90_658 ();
 FILLCELL_X2 FILLER_90_662 ();
 FILLCELL_X16 FILLER_90_673 ();
 FILLCELL_X8 FILLER_90_702 ();
 FILLCELL_X4 FILLER_90_710 ();
 FILLCELL_X4 FILLER_90_725 ();
 FILLCELL_X2 FILLER_90_729 ();
 FILLCELL_X1 FILLER_90_731 ();
 FILLCELL_X2 FILLER_90_750 ();
 FILLCELL_X1 FILLER_90_752 ();
 FILLCELL_X4 FILLER_90_767 ();
 FILLCELL_X2 FILLER_90_771 ();
 FILLCELL_X1 FILLER_90_776 ();
 FILLCELL_X2 FILLER_90_780 ();
 FILLCELL_X1 FILLER_90_793 ();
 FILLCELL_X2 FILLER_90_800 ();
 FILLCELL_X1 FILLER_90_817 ();
 FILLCELL_X4 FILLER_90_829 ();
 FILLCELL_X4 FILLER_90_836 ();
 FILLCELL_X1 FILLER_90_840 ();
 FILLCELL_X4 FILLER_90_857 ();
 FILLCELL_X2 FILLER_90_861 ();
 FILLCELL_X1 FILLER_90_863 ();
 FILLCELL_X16 FILLER_90_867 ();
 FILLCELL_X1 FILLER_90_883 ();
 FILLCELL_X8 FILLER_90_888 ();
 FILLCELL_X2 FILLER_90_896 ();
 FILLCELL_X1 FILLER_90_898 ();
 FILLCELL_X4 FILLER_90_911 ();
 FILLCELL_X2 FILLER_90_915 ();
 FILLCELL_X2 FILLER_90_930 ();
 FILLCELL_X2 FILLER_90_939 ();
 FILLCELL_X1 FILLER_90_941 ();
 FILLCELL_X16 FILLER_90_953 ();
 FILLCELL_X4 FILLER_90_980 ();
 FILLCELL_X2 FILLER_90_984 ();
 FILLCELL_X1 FILLER_90_986 ();
 FILLCELL_X2 FILLER_90_1008 ();
 FILLCELL_X1 FILLER_90_1010 ();
 FILLCELL_X8 FILLER_90_1022 ();
 FILLCELL_X1 FILLER_90_1030 ();
 FILLCELL_X1 FILLER_90_1035 ();
 FILLCELL_X1 FILLER_90_1038 ();
 FILLCELL_X2 FILLER_90_1045 ();
 FILLCELL_X1 FILLER_90_1064 ();
 FILLCELL_X4 FILLER_90_1069 ();
 FILLCELL_X2 FILLER_90_1080 ();
 FILLCELL_X1 FILLER_90_1082 ();
 FILLCELL_X4 FILLER_90_1090 ();
 FILLCELL_X1 FILLER_90_1094 ();
 FILLCELL_X4 FILLER_90_1105 ();
 FILLCELL_X4 FILLER_90_1113 ();
 FILLCELL_X1 FILLER_90_1120 ();
 FILLCELL_X1 FILLER_90_1124 ();
 FILLCELL_X2 FILLER_90_1130 ();
 FILLCELL_X1 FILLER_90_1132 ();
 FILLCELL_X2 FILLER_90_1139 ();
 FILLCELL_X2 FILLER_90_1165 ();
 FILLCELL_X8 FILLER_90_1171 ();
 FILLCELL_X2 FILLER_90_1224 ();
 FILLCELL_X1 FILLER_90_1228 ();
 FILLCELL_X4 FILLER_90_1242 ();
 FILLCELL_X1 FILLER_90_1246 ();
 FILLCELL_X2 FILLER_90_1250 ();
 FILLCELL_X2 FILLER_91_1 ();
 FILLCELL_X1 FILLER_91_3 ();
 FILLCELL_X4 FILLER_91_24 ();
 FILLCELL_X4 FILLER_91_35 ();
 FILLCELL_X2 FILLER_91_39 ();
 FILLCELL_X8 FILLER_91_48 ();
 FILLCELL_X2 FILLER_91_56 ();
 FILLCELL_X1 FILLER_91_58 ();
 FILLCELL_X4 FILLER_91_66 ();
 FILLCELL_X8 FILLER_91_77 ();
 FILLCELL_X4 FILLER_91_85 ();
 FILLCELL_X1 FILLER_91_89 ();
 FILLCELL_X1 FILLER_91_97 ();
 FILLCELL_X1 FILLER_91_105 ();
 FILLCELL_X16 FILLER_91_113 ();
 FILLCELL_X1 FILLER_91_129 ();
 FILLCELL_X4 FILLER_91_137 ();
 FILLCELL_X1 FILLER_91_148 ();
 FILLCELL_X2 FILLER_91_186 ();
 FILLCELL_X16 FILLER_91_195 ();
 FILLCELL_X4 FILLER_91_211 ();
 FILLCELL_X1 FILLER_91_219 ();
 FILLCELL_X4 FILLER_91_230 ();
 FILLCELL_X4 FILLER_91_238 ();
 FILLCELL_X1 FILLER_91_242 ();
 FILLCELL_X4 FILLER_91_246 ();
 FILLCELL_X1 FILLER_91_250 ();
 FILLCELL_X4 FILLER_91_281 ();
 FILLCELL_X1 FILLER_91_285 ();
 FILLCELL_X1 FILLER_91_302 ();
 FILLCELL_X2 FILLER_91_307 ();
 FILLCELL_X16 FILLER_91_316 ();
 FILLCELL_X8 FILLER_91_332 ();
 FILLCELL_X1 FILLER_91_340 ();
 FILLCELL_X4 FILLER_91_372 ();
 FILLCELL_X2 FILLER_91_376 ();
 FILLCELL_X8 FILLER_91_394 ();
 FILLCELL_X2 FILLER_91_402 ();
 FILLCELL_X1 FILLER_91_404 ();
 FILLCELL_X4 FILLER_91_409 ();
 FILLCELL_X1 FILLER_91_413 ();
 FILLCELL_X1 FILLER_91_421 ();
 FILLCELL_X1 FILLER_91_429 ();
 FILLCELL_X2 FILLER_91_437 ();
 FILLCELL_X4 FILLER_91_446 ();
 FILLCELL_X1 FILLER_91_450 ();
 FILLCELL_X2 FILLER_91_461 ();
 FILLCELL_X8 FILLER_91_472 ();
 FILLCELL_X1 FILLER_91_480 ();
 FILLCELL_X4 FILLER_91_486 ();
 FILLCELL_X2 FILLER_91_490 ();
 FILLCELL_X8 FILLER_91_499 ();
 FILLCELL_X2 FILLER_91_507 ();
 FILLCELL_X1 FILLER_91_509 ();
 FILLCELL_X4 FILLER_91_523 ();
 FILLCELL_X2 FILLER_91_527 ();
 FILLCELL_X1 FILLER_91_571 ();
 FILLCELL_X1 FILLER_91_592 ();
 FILLCELL_X2 FILLER_91_607 ();
 FILLCELL_X8 FILLER_91_616 ();
 FILLCELL_X1 FILLER_91_624 ();
 FILLCELL_X2 FILLER_91_636 ();
 FILLCELL_X1 FILLER_91_638 ();
 FILLCELL_X8 FILLER_91_654 ();
 FILLCELL_X2 FILLER_91_662 ();
 FILLCELL_X1 FILLER_91_676 ();
 FILLCELL_X4 FILLER_91_690 ();
 FILLCELL_X2 FILLER_91_694 ();
 FILLCELL_X1 FILLER_91_696 ();
 FILLCELL_X8 FILLER_91_702 ();
 FILLCELL_X4 FILLER_91_710 ();
 FILLCELL_X2 FILLER_91_714 ();
 FILLCELL_X32 FILLER_91_723 ();
 FILLCELL_X16 FILLER_91_755 ();
 FILLCELL_X2 FILLER_91_771 ();
 FILLCELL_X1 FILLER_91_773 ();
 FILLCELL_X8 FILLER_91_781 ();
 FILLCELL_X2 FILLER_91_789 ();
 FILLCELL_X1 FILLER_91_791 ();
 FILLCELL_X8 FILLER_91_800 ();
 FILLCELL_X8 FILLER_91_816 ();
 FILLCELL_X2 FILLER_91_824 ();
 FILLCELL_X1 FILLER_91_826 ();
 FILLCELL_X8 FILLER_91_848 ();
 FILLCELL_X2 FILLER_91_856 ();
 FILLCELL_X1 FILLER_91_858 ();
 FILLCELL_X4 FILLER_91_869 ();
 FILLCELL_X2 FILLER_91_873 ();
 FILLCELL_X8 FILLER_91_885 ();
 FILLCELL_X4 FILLER_91_893 ();
 FILLCELL_X2 FILLER_91_897 ();
 FILLCELL_X8 FILLER_91_902 ();
 FILLCELL_X1 FILLER_91_910 ();
 FILLCELL_X1 FILLER_91_924 ();
 FILLCELL_X4 FILLER_91_972 ();
 FILLCELL_X1 FILLER_91_976 ();
 FILLCELL_X1 FILLER_91_984 ();
 FILLCELL_X4 FILLER_91_1012 ();
 FILLCELL_X2 FILLER_91_1016 ();
 FILLCELL_X1 FILLER_91_1018 ();
 FILLCELL_X4 FILLER_91_1023 ();
 FILLCELL_X2 FILLER_91_1027 ();
 FILLCELL_X1 FILLER_91_1038 ();
 FILLCELL_X2 FILLER_91_1043 ();
 FILLCELL_X1 FILLER_91_1045 ();
 FILLCELL_X8 FILLER_91_1052 ();
 FILLCELL_X1 FILLER_91_1060 ();
 FILLCELL_X8 FILLER_91_1065 ();
 FILLCELL_X4 FILLER_91_1073 ();
 FILLCELL_X2 FILLER_91_1077 ();
 FILLCELL_X4 FILLER_91_1097 ();
 FILLCELL_X4 FILLER_91_1109 ();
 FILLCELL_X2 FILLER_91_1113 ();
 FILLCELL_X1 FILLER_91_1115 ();
 FILLCELL_X4 FILLER_91_1128 ();
 FILLCELL_X1 FILLER_91_1132 ();
 FILLCELL_X4 FILLER_91_1169 ();
 FILLCELL_X2 FILLER_91_1173 ();
 FILLCELL_X1 FILLER_91_1175 ();
 FILLCELL_X8 FILLER_91_1205 ();
 FILLCELL_X4 FILLER_91_1213 ();
 FILLCELL_X2 FILLER_91_1217 ();
 FILLCELL_X2 FILLER_91_1236 ();
 FILLCELL_X8 FILLER_92_1 ();
 FILLCELL_X4 FILLER_92_43 ();
 FILLCELL_X4 FILLER_92_67 ();
 FILLCELL_X4 FILLER_92_98 ();
 FILLCELL_X1 FILLER_92_102 ();
 FILLCELL_X2 FILLER_92_110 ();
 FILLCELL_X1 FILLER_92_112 ();
 FILLCELL_X2 FILLER_92_154 ();
 FILLCELL_X1 FILLER_92_156 ();
 FILLCELL_X2 FILLER_92_177 ();
 FILLCELL_X1 FILLER_92_179 ();
 FILLCELL_X2 FILLER_92_224 ();
 FILLCELL_X1 FILLER_92_226 ();
 FILLCELL_X1 FILLER_92_247 ();
 FILLCELL_X2 FILLER_92_275 ();
 FILLCELL_X1 FILLER_92_322 ();
 FILLCELL_X4 FILLER_92_331 ();
 FILLCELL_X1 FILLER_92_382 ();
 FILLCELL_X4 FILLER_92_397 ();
 FILLCELL_X2 FILLER_92_421 ();
 FILLCELL_X4 FILLER_92_446 ();
 FILLCELL_X2 FILLER_92_450 ();
 FILLCELL_X2 FILLER_92_456 ();
 FILLCELL_X2 FILLER_92_475 ();
 FILLCELL_X2 FILLER_92_490 ();
 FILLCELL_X1 FILLER_92_492 ();
 FILLCELL_X8 FILLER_92_506 ();
 FILLCELL_X4 FILLER_92_514 ();
 FILLCELL_X4 FILLER_92_525 ();
 FILLCELL_X2 FILLER_92_529 ();
 FILLCELL_X1 FILLER_92_531 ();
 FILLCELL_X16 FILLER_92_579 ();
 FILLCELL_X4 FILLER_92_595 ();
 FILLCELL_X2 FILLER_92_619 ();
 FILLCELL_X2 FILLER_92_641 ();
 FILLCELL_X1 FILLER_92_653 ();
 FILLCELL_X1 FILLER_92_668 ();
 FILLCELL_X1 FILLER_92_679 ();
 FILLCELL_X2 FILLER_92_685 ();
 FILLCELL_X1 FILLER_92_687 ();
 FILLCELL_X2 FILLER_92_697 ();
 FILLCELL_X1 FILLER_92_699 ();
 FILLCELL_X16 FILLER_92_721 ();
 FILLCELL_X8 FILLER_92_737 ();
 FILLCELL_X4 FILLER_92_745 ();
 FILLCELL_X4 FILLER_92_767 ();
 FILLCELL_X4 FILLER_92_789 ();
 FILLCELL_X2 FILLER_92_804 ();
 FILLCELL_X1 FILLER_92_806 ();
 FILLCELL_X2 FILLER_92_840 ();
 FILLCELL_X1 FILLER_92_842 ();
 FILLCELL_X2 FILLER_92_879 ();
 FILLCELL_X1 FILLER_92_881 ();
 FILLCELL_X4 FILLER_92_913 ();
 FILLCELL_X2 FILLER_92_917 ();
 FILLCELL_X1 FILLER_92_927 ();
 FILLCELL_X16 FILLER_92_935 ();
 FILLCELL_X4 FILLER_92_951 ();
 FILLCELL_X2 FILLER_92_955 ();
 FILLCELL_X4 FILLER_92_971 ();
 FILLCELL_X1 FILLER_92_984 ();
 FILLCELL_X8 FILLER_92_996 ();
 FILLCELL_X2 FILLER_92_1004 ();
 FILLCELL_X1 FILLER_92_1006 ();
 FILLCELL_X1 FILLER_92_1031 ();
 FILLCELL_X8 FILLER_92_1045 ();
 FILLCELL_X2 FILLER_92_1053 ();
 FILLCELL_X4 FILLER_92_1076 ();
 FILLCELL_X2 FILLER_92_1099 ();
 FILLCELL_X4 FILLER_92_1116 ();
 FILLCELL_X2 FILLER_92_1120 ();
 FILLCELL_X1 FILLER_92_1122 ();
 FILLCELL_X1 FILLER_92_1127 ();
 FILLCELL_X8 FILLER_92_1133 ();
 FILLCELL_X2 FILLER_92_1141 ();
 FILLCELL_X1 FILLER_92_1143 ();
 FILLCELL_X8 FILLER_92_1161 ();
 FILLCELL_X2 FILLER_92_1169 ();
 FILLCELL_X1 FILLER_92_1175 ();
 FILLCELL_X2 FILLER_92_1180 ();
 FILLCELL_X16 FILLER_92_1196 ();
 FILLCELL_X2 FILLER_92_1212 ();
 FILLCELL_X4 FILLER_92_1227 ();
 FILLCELL_X1 FILLER_92_1245 ();
 FILLCELL_X2 FILLER_92_1252 ();
 FILLCELL_X1 FILLER_92_1254 ();
 FILLCELL_X16 FILLER_93_1 ();
 FILLCELL_X2 FILLER_93_17 ();
 FILLCELL_X4 FILLER_93_26 ();
 FILLCELL_X2 FILLER_93_30 ();
 FILLCELL_X1 FILLER_93_32 ();
 FILLCELL_X4 FILLER_93_67 ();
 FILLCELL_X2 FILLER_93_98 ();
 FILLCELL_X1 FILLER_93_100 ();
 FILLCELL_X1 FILLER_93_108 ();
 FILLCELL_X1 FILLER_93_136 ();
 FILLCELL_X8 FILLER_93_151 ();
 FILLCELL_X2 FILLER_93_159 ();
 FILLCELL_X1 FILLER_93_161 ();
 FILLCELL_X16 FILLER_93_169 ();
 FILLCELL_X1 FILLER_93_185 ();
 FILLCELL_X2 FILLER_93_200 ();
 FILLCELL_X1 FILLER_93_222 ();
 FILLCELL_X8 FILLER_93_249 ();
 FILLCELL_X2 FILLER_93_257 ();
 FILLCELL_X1 FILLER_93_259 ();
 FILLCELL_X2 FILLER_93_309 ();
 FILLCELL_X1 FILLER_93_326 ();
 FILLCELL_X8 FILLER_93_337 ();
 FILLCELL_X2 FILLER_93_345 ();
 FILLCELL_X4 FILLER_93_351 ();
 FILLCELL_X2 FILLER_93_355 ();
 FILLCELL_X4 FILLER_93_360 ();
 FILLCELL_X8 FILLER_93_374 ();
 FILLCELL_X2 FILLER_93_382 ();
 FILLCELL_X1 FILLER_93_384 ();
 FILLCELL_X2 FILLER_93_392 ();
 FILLCELL_X1 FILLER_93_394 ();
 FILLCELL_X2 FILLER_93_402 ();
 FILLCELL_X8 FILLER_93_414 ();
 FILLCELL_X4 FILLER_93_422 ();
 FILLCELL_X2 FILLER_93_426 ();
 FILLCELL_X1 FILLER_93_428 ();
 FILLCELL_X4 FILLER_93_433 ();
 FILLCELL_X2 FILLER_93_437 ();
 FILLCELL_X4 FILLER_93_446 ();
 FILLCELL_X1 FILLER_93_450 ();
 FILLCELL_X8 FILLER_93_454 ();
 FILLCELL_X2 FILLER_93_465 ();
 FILLCELL_X1 FILLER_93_467 ();
 FILLCELL_X4 FILLER_93_475 ();
 FILLCELL_X2 FILLER_93_479 ();
 FILLCELL_X8 FILLER_93_553 ();
 FILLCELL_X8 FILLER_93_595 ();
 FILLCELL_X16 FILLER_93_610 ();
 FILLCELL_X4 FILLER_93_626 ();
 FILLCELL_X1 FILLER_93_630 ();
 FILLCELL_X2 FILLER_93_644 ();
 FILLCELL_X1 FILLER_93_646 ();
 FILLCELL_X8 FILLER_93_649 ();
 FILLCELL_X4 FILLER_93_657 ();
 FILLCELL_X2 FILLER_93_661 ();
 FILLCELL_X1 FILLER_93_663 ();
 FILLCELL_X1 FILLER_93_676 ();
 FILLCELL_X2 FILLER_93_691 ();
 FILLCELL_X1 FILLER_93_700 ();
 FILLCELL_X1 FILLER_93_704 ();
 FILLCELL_X1 FILLER_93_709 ();
 FILLCELL_X1 FILLER_93_724 ();
 FILLCELL_X16 FILLER_93_738 ();
 FILLCELL_X4 FILLER_93_754 ();
 FILLCELL_X2 FILLER_93_758 ();
 FILLCELL_X1 FILLER_93_767 ();
 FILLCELL_X1 FILLER_93_777 ();
 FILLCELL_X8 FILLER_93_802 ();
 FILLCELL_X2 FILLER_93_810 ();
 FILLCELL_X1 FILLER_93_815 ();
 FILLCELL_X2 FILLER_93_825 ();
 FILLCELL_X2 FILLER_93_837 ();
 FILLCELL_X4 FILLER_93_841 ();
 FILLCELL_X4 FILLER_93_871 ();
 FILLCELL_X2 FILLER_93_875 ();
 FILLCELL_X4 FILLER_93_888 ();
 FILLCELL_X2 FILLER_93_892 ();
 FILLCELL_X8 FILLER_93_908 ();
 FILLCELL_X4 FILLER_93_916 ();
 FILLCELL_X1 FILLER_93_920 ();
 FILLCELL_X1 FILLER_93_924 ();
 FILLCELL_X2 FILLER_93_952 ();
 FILLCELL_X2 FILLER_93_961 ();
 FILLCELL_X4 FILLER_93_970 ();
 FILLCELL_X4 FILLER_93_991 ();
 FILLCELL_X8 FILLER_93_1002 ();
 FILLCELL_X4 FILLER_93_1010 ();
 FILLCELL_X1 FILLER_93_1014 ();
 FILLCELL_X1 FILLER_93_1034 ();
 FILLCELL_X8 FILLER_93_1039 ();
 FILLCELL_X2 FILLER_93_1047 ();
 FILLCELL_X4 FILLER_93_1062 ();
 FILLCELL_X1 FILLER_93_1066 ();
 FILLCELL_X4 FILLER_93_1070 ();
 FILLCELL_X1 FILLER_93_1095 ();
 FILLCELL_X4 FILLER_93_1109 ();
 FILLCELL_X2 FILLER_93_1113 ();
 FILLCELL_X1 FILLER_93_1115 ();
 FILLCELL_X1 FILLER_93_1133 ();
 FILLCELL_X1 FILLER_93_1160 ();
 FILLCELL_X2 FILLER_93_1180 ();
 FILLCELL_X1 FILLER_93_1182 ();
 FILLCELL_X4 FILLER_93_1192 ();
 FILLCELL_X1 FILLER_93_1196 ();
 FILLCELL_X1 FILLER_93_1208 ();
 FILLCELL_X4 FILLER_93_1233 ();
 FILLCELL_X1 FILLER_93_1237 ();
 FILLCELL_X4 FILLER_94_28 ();
 FILLCELL_X1 FILLER_94_32 ();
 FILLCELL_X8 FILLER_94_40 ();
 FILLCELL_X2 FILLER_94_48 ();
 FILLCELL_X1 FILLER_94_50 ();
 FILLCELL_X4 FILLER_94_76 ();
 FILLCELL_X1 FILLER_94_80 ();
 FILLCELL_X4 FILLER_94_88 ();
 FILLCELL_X1 FILLER_94_92 ();
 FILLCELL_X16 FILLER_94_107 ();
 FILLCELL_X8 FILLER_94_150 ();
 FILLCELL_X1 FILLER_94_165 ();
 FILLCELL_X1 FILLER_94_186 ();
 FILLCELL_X16 FILLER_94_201 ();
 FILLCELL_X1 FILLER_94_217 ();
 FILLCELL_X4 FILLER_94_226 ();
 FILLCELL_X2 FILLER_94_230 ();
 FILLCELL_X1 FILLER_94_232 ();
 FILLCELL_X4 FILLER_94_237 ();
 FILLCELL_X1 FILLER_94_241 ();
 FILLCELL_X4 FILLER_94_250 ();
 FILLCELL_X1 FILLER_94_261 ();
 FILLCELL_X2 FILLER_94_282 ();
 FILLCELL_X1 FILLER_94_294 ();
 FILLCELL_X1 FILLER_94_309 ();
 FILLCELL_X2 FILLER_94_317 ();
 FILLCELL_X2 FILLER_94_344 ();
 FILLCELL_X4 FILLER_94_366 ();
 FILLCELL_X2 FILLER_94_370 ();
 FILLCELL_X1 FILLER_94_398 ();
 FILLCELL_X2 FILLER_94_427 ();
 FILLCELL_X1 FILLER_94_429 ();
 FILLCELL_X2 FILLER_94_434 ();
 FILLCELL_X8 FILLER_94_453 ();
 FILLCELL_X4 FILLER_94_461 ();
 FILLCELL_X1 FILLER_94_485 ();
 FILLCELL_X4 FILLER_94_534 ();
 FILLCELL_X1 FILLER_94_538 ();
 FILLCELL_X16 FILLER_94_543 ();
 FILLCELL_X4 FILLER_94_559 ();
 FILLCELL_X1 FILLER_94_563 ();
 FILLCELL_X2 FILLER_94_619 ();
 FILLCELL_X1 FILLER_94_632 ();
 FILLCELL_X4 FILLER_94_646 ();
 FILLCELL_X2 FILLER_94_650 ();
 FILLCELL_X1 FILLER_94_652 ();
 FILLCELL_X1 FILLER_94_675 ();
 FILLCELL_X1 FILLER_94_679 ();
 FILLCELL_X2 FILLER_94_692 ();
 FILLCELL_X2 FILLER_94_702 ();
 FILLCELL_X4 FILLER_94_724 ();
 FILLCELL_X1 FILLER_94_733 ();
 FILLCELL_X1 FILLER_94_738 ();
 FILLCELL_X2 FILLER_94_743 ();
 FILLCELL_X1 FILLER_94_749 ();
 FILLCELL_X4 FILLER_94_754 ();
 FILLCELL_X2 FILLER_94_758 ();
 FILLCELL_X4 FILLER_94_774 ();
 FILLCELL_X2 FILLER_94_778 ();
 FILLCELL_X16 FILLER_94_783 ();
 FILLCELL_X4 FILLER_94_799 ();
 FILLCELL_X1 FILLER_94_803 ();
 FILLCELL_X8 FILLER_94_806 ();
 FILLCELL_X1 FILLER_94_814 ();
 FILLCELL_X8 FILLER_94_821 ();
 FILLCELL_X4 FILLER_94_829 ();
 FILLCELL_X1 FILLER_94_833 ();
 FILLCELL_X2 FILLER_94_847 ();
 FILLCELL_X1 FILLER_94_849 ();
 FILLCELL_X4 FILLER_94_868 ();
 FILLCELL_X2 FILLER_94_872 ();
 FILLCELL_X1 FILLER_94_900 ();
 FILLCELL_X2 FILLER_94_904 ();
 FILLCELL_X1 FILLER_94_906 ();
 FILLCELL_X2 FILLER_94_909 ();
 FILLCELL_X2 FILLER_94_923 ();
 FILLCELL_X8 FILLER_94_928 ();
 FILLCELL_X4 FILLER_94_936 ();
 FILLCELL_X1 FILLER_94_940 ();
 FILLCELL_X1 FILLER_94_948 ();
 FILLCELL_X2 FILLER_94_963 ();
 FILLCELL_X2 FILLER_94_987 ();
 FILLCELL_X2 FILLER_94_1011 ();
 FILLCELL_X1 FILLER_94_1013 ();
 FILLCELL_X8 FILLER_94_1022 ();
 FILLCELL_X4 FILLER_94_1030 ();
 FILLCELL_X4 FILLER_94_1042 ();
 FILLCELL_X8 FILLER_94_1055 ();
 FILLCELL_X2 FILLER_94_1063 ();
 FILLCELL_X8 FILLER_94_1106 ();
 FILLCELL_X2 FILLER_94_1114 ();
 FILLCELL_X1 FILLER_94_1116 ();
 FILLCELL_X8 FILLER_94_1123 ();
 FILLCELL_X1 FILLER_94_1137 ();
 FILLCELL_X2 FILLER_94_1142 ();
 FILLCELL_X1 FILLER_94_1144 ();
 FILLCELL_X8 FILLER_94_1149 ();
 FILLCELL_X2 FILLER_94_1157 ();
 FILLCELL_X4 FILLER_94_1169 ();
 FILLCELL_X1 FILLER_94_1173 ();
 FILLCELL_X4 FILLER_94_1183 ();
 FILLCELL_X1 FILLER_94_1187 ();
 FILLCELL_X1 FILLER_94_1208 ();
 FILLCELL_X2 FILLER_94_1217 ();
 FILLCELL_X1 FILLER_94_1219 ();
 FILLCELL_X2 FILLER_94_1222 ();
 FILLCELL_X2 FILLER_94_1229 ();
 FILLCELL_X4 FILLER_94_1245 ();
 FILLCELL_X2 FILLER_94_1249 ();
 FILLCELL_X1 FILLER_94_1251 ();
 FILLCELL_X16 FILLER_95_1 ();
 FILLCELL_X2 FILLER_95_17 ();
 FILLCELL_X4 FILLER_95_39 ();
 FILLCELL_X2 FILLER_95_43 ();
 FILLCELL_X1 FILLER_95_45 ();
 FILLCELL_X4 FILLER_95_53 ();
 FILLCELL_X1 FILLER_95_57 ();
 FILLCELL_X2 FILLER_95_61 ();
 FILLCELL_X1 FILLER_95_70 ();
 FILLCELL_X1 FILLER_95_78 ();
 FILLCELL_X2 FILLER_95_113 ();
 FILLCELL_X1 FILLER_95_115 ();
 FILLCELL_X16 FILLER_95_127 ();
 FILLCELL_X1 FILLER_95_143 ();
 FILLCELL_X8 FILLER_95_171 ();
 FILLCELL_X4 FILLER_95_179 ();
 FILLCELL_X1 FILLER_95_183 ();
 FILLCELL_X1 FILLER_95_198 ();
 FILLCELL_X1 FILLER_95_245 ();
 FILLCELL_X1 FILLER_95_273 ();
 FILLCELL_X4 FILLER_95_299 ();
 FILLCELL_X1 FILLER_95_303 ();
 FILLCELL_X4 FILLER_95_307 ();
 FILLCELL_X2 FILLER_95_311 ();
 FILLCELL_X8 FILLER_95_336 ();
 FILLCELL_X2 FILLER_95_344 ();
 FILLCELL_X1 FILLER_95_346 ();
 FILLCELL_X1 FILLER_95_351 ();
 FILLCELL_X4 FILLER_95_356 ();
 FILLCELL_X1 FILLER_95_360 ();
 FILLCELL_X16 FILLER_95_364 ();
 FILLCELL_X2 FILLER_95_388 ();
 FILLCELL_X8 FILLER_95_400 ();
 FILLCELL_X8 FILLER_95_415 ();
 FILLCELL_X2 FILLER_95_423 ();
 FILLCELL_X1 FILLER_95_425 ();
 FILLCELL_X2 FILLER_95_453 ();
 FILLCELL_X4 FILLER_95_478 ();
 FILLCELL_X1 FILLER_95_482 ();
 FILLCELL_X2 FILLER_95_503 ();
 FILLCELL_X1 FILLER_95_505 ();
 FILLCELL_X8 FILLER_95_540 ();
 FILLCELL_X1 FILLER_95_548 ();
 FILLCELL_X1 FILLER_95_556 ();
 FILLCELL_X2 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_586 ();
 FILLCELL_X1 FILLER_95_618 ();
 FILLCELL_X8 FILLER_95_636 ();
 FILLCELL_X2 FILLER_95_644 ();
 FILLCELL_X1 FILLER_95_646 ();
 FILLCELL_X8 FILLER_95_656 ();
 FILLCELL_X4 FILLER_95_664 ();
 FILLCELL_X1 FILLER_95_680 ();
 FILLCELL_X8 FILLER_95_689 ();
 FILLCELL_X2 FILLER_95_697 ();
 FILLCELL_X1 FILLER_95_699 ();
 FILLCELL_X4 FILLER_95_710 ();
 FILLCELL_X2 FILLER_95_714 ();
 FILLCELL_X1 FILLER_95_716 ();
 FILLCELL_X8 FILLER_95_729 ();
 FILLCELL_X2 FILLER_95_737 ();
 FILLCELL_X1 FILLER_95_739 ();
 FILLCELL_X2 FILLER_95_755 ();
 FILLCELL_X1 FILLER_95_757 ();
 FILLCELL_X1 FILLER_95_770 ();
 FILLCELL_X8 FILLER_95_786 ();
 FILLCELL_X2 FILLER_95_825 ();
 FILLCELL_X4 FILLER_95_843 ();
 FILLCELL_X1 FILLER_95_847 ();
 FILLCELL_X4 FILLER_95_876 ();
 FILLCELL_X2 FILLER_95_887 ();
 FILLCELL_X2 FILLER_95_895 ();
 FILLCELL_X1 FILLER_95_897 ();
 FILLCELL_X16 FILLER_95_913 ();
 FILLCELL_X8 FILLER_95_929 ();
 FILLCELL_X2 FILLER_95_937 ();
 FILLCELL_X1 FILLER_95_973 ();
 FILLCELL_X4 FILLER_95_977 ();
 FILLCELL_X1 FILLER_95_981 ();
 FILLCELL_X4 FILLER_95_999 ();
 FILLCELL_X1 FILLER_95_1003 ();
 FILLCELL_X8 FILLER_95_1025 ();
 FILLCELL_X4 FILLER_95_1033 ();
 FILLCELL_X1 FILLER_95_1037 ();
 FILLCELL_X1 FILLER_95_1053 ();
 FILLCELL_X8 FILLER_95_1080 ();
 FILLCELL_X2 FILLER_95_1088 ();
 FILLCELL_X8 FILLER_95_1094 ();
 FILLCELL_X2 FILLER_95_1102 ();
 FILLCELL_X4 FILLER_95_1147 ();
 FILLCELL_X8 FILLER_95_1154 ();
 FILLCELL_X2 FILLER_95_1162 ();
 FILLCELL_X1 FILLER_95_1164 ();
 FILLCELL_X1 FILLER_95_1167 ();
 FILLCELL_X2 FILLER_95_1175 ();
 FILLCELL_X1 FILLER_95_1203 ();
 FILLCELL_X2 FILLER_95_1221 ();
 FILLCELL_X2 FILLER_95_1229 ();
 FILLCELL_X1 FILLER_95_1238 ();
 FILLCELL_X2 FILLER_95_1253 ();
 FILLCELL_X8 FILLER_96_1 ();
 FILLCELL_X4 FILLER_96_9 ();
 FILLCELL_X2 FILLER_96_13 ();
 FILLCELL_X1 FILLER_96_15 ();
 FILLCELL_X2 FILLER_96_30 ();
 FILLCELL_X1 FILLER_96_32 ();
 FILLCELL_X16 FILLER_96_40 ();
 FILLCELL_X4 FILLER_96_56 ();
 FILLCELL_X2 FILLER_96_87 ();
 FILLCELL_X1 FILLER_96_103 ();
 FILLCELL_X8 FILLER_96_111 ();
 FILLCELL_X2 FILLER_96_123 ();
 FILLCELL_X1 FILLER_96_125 ();
 FILLCELL_X16 FILLER_96_158 ();
 FILLCELL_X4 FILLER_96_174 ();
 FILLCELL_X8 FILLER_96_198 ();
 FILLCELL_X4 FILLER_96_206 ();
 FILLCELL_X1 FILLER_96_210 ();
 FILLCELL_X8 FILLER_96_225 ();
 FILLCELL_X1 FILLER_96_237 ();
 FILLCELL_X1 FILLER_96_242 ();
 FILLCELL_X1 FILLER_96_246 ();
 FILLCELL_X2 FILLER_96_254 ();
 FILLCELL_X2 FILLER_96_261 ();
 FILLCELL_X1 FILLER_96_263 ();
 FILLCELL_X2 FILLER_96_284 ();
 FILLCELL_X1 FILLER_96_286 ();
 FILLCELL_X2 FILLER_96_307 ();
 FILLCELL_X1 FILLER_96_309 ();
 FILLCELL_X8 FILLER_96_330 ();
 FILLCELL_X1 FILLER_96_338 ();
 FILLCELL_X2 FILLER_96_362 ();
 FILLCELL_X1 FILLER_96_374 ();
 FILLCELL_X2 FILLER_96_379 ();
 FILLCELL_X2 FILLER_96_401 ();
 FILLCELL_X2 FILLER_96_410 ();
 FILLCELL_X1 FILLER_96_412 ();
 FILLCELL_X8 FILLER_96_420 ();
 FILLCELL_X1 FILLER_96_428 ();
 FILLCELL_X8 FILLER_96_433 ();
 FILLCELL_X1 FILLER_96_441 ();
 FILLCELL_X8 FILLER_96_452 ();
 FILLCELL_X4 FILLER_96_460 ();
 FILLCELL_X1 FILLER_96_464 ();
 FILLCELL_X2 FILLER_96_479 ();
 FILLCELL_X1 FILLER_96_481 ();
 FILLCELL_X4 FILLER_96_489 ();
 FILLCELL_X2 FILLER_96_500 ();
 FILLCELL_X1 FILLER_96_502 ();
 FILLCELL_X2 FILLER_96_510 ();
 FILLCELL_X4 FILLER_96_519 ();
 FILLCELL_X4 FILLER_96_530 ();
 FILLCELL_X4 FILLER_96_541 ();
 FILLCELL_X2 FILLER_96_545 ();
 FILLCELL_X8 FILLER_96_561 ();
 FILLCELL_X4 FILLER_96_569 ();
 FILLCELL_X1 FILLER_96_573 ();
 FILLCELL_X8 FILLER_96_581 ();
 FILLCELL_X1 FILLER_96_589 ();
 FILLCELL_X8 FILLER_96_617 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X16 FILLER_96_632 ();
 FILLCELL_X1 FILLER_96_705 ();
 FILLCELL_X2 FILLER_96_719 ();
 FILLCELL_X2 FILLER_96_726 ();
 FILLCELL_X1 FILLER_96_732 ();
 FILLCELL_X2 FILLER_96_738 ();
 FILLCELL_X1 FILLER_96_744 ();
 FILLCELL_X2 FILLER_96_749 ();
 FILLCELL_X32 FILLER_96_755 ();
 FILLCELL_X8 FILLER_96_787 ();
 FILLCELL_X1 FILLER_96_799 ();
 FILLCELL_X4 FILLER_96_815 ();
 FILLCELL_X1 FILLER_96_823 ();
 FILLCELL_X4 FILLER_96_840 ();
 FILLCELL_X2 FILLER_96_844 ();
 FILLCELL_X1 FILLER_96_846 ();
 FILLCELL_X1 FILLER_96_862 ();
 FILLCELL_X2 FILLER_96_870 ();
 FILLCELL_X1 FILLER_96_872 ();
 FILLCELL_X8 FILLER_96_878 ();
 FILLCELL_X2 FILLER_96_886 ();
 FILLCELL_X1 FILLER_96_888 ();
 FILLCELL_X8 FILLER_96_894 ();
 FILLCELL_X2 FILLER_96_902 ();
 FILLCELL_X1 FILLER_96_904 ();
 FILLCELL_X4 FILLER_96_908 ();
 FILLCELL_X2 FILLER_96_912 ();
 FILLCELL_X2 FILLER_96_923 ();
 FILLCELL_X4 FILLER_96_930 ();
 FILLCELL_X1 FILLER_96_934 ();
 FILLCELL_X1 FILLER_96_944 ();
 FILLCELL_X2 FILLER_96_948 ();
 FILLCELL_X1 FILLER_96_950 ();
 FILLCELL_X8 FILLER_96_958 ();
 FILLCELL_X2 FILLER_96_966 ();
 FILLCELL_X4 FILLER_96_985 ();
 FILLCELL_X1 FILLER_96_989 ();
 FILLCELL_X16 FILLER_96_1007 ();
 FILLCELL_X4 FILLER_96_1023 ();
 FILLCELL_X2 FILLER_96_1027 ();
 FILLCELL_X4 FILLER_96_1051 ();
 FILLCELL_X2 FILLER_96_1055 ();
 FILLCELL_X1 FILLER_96_1064 ();
 FILLCELL_X16 FILLER_96_1067 ();
 FILLCELL_X2 FILLER_96_1083 ();
 FILLCELL_X1 FILLER_96_1085 ();
 FILLCELL_X4 FILLER_96_1110 ();
 FILLCELL_X4 FILLER_96_1117 ();
 FILLCELL_X2 FILLER_96_1125 ();
 FILLCELL_X1 FILLER_96_1127 ();
 FILLCELL_X2 FILLER_96_1144 ();
 FILLCELL_X1 FILLER_96_1146 ();
 FILLCELL_X8 FILLER_96_1181 ();
 FILLCELL_X2 FILLER_96_1206 ();
 FILLCELL_X4 FILLER_96_1213 ();
 FILLCELL_X1 FILLER_96_1228 ();
 FILLCELL_X4 FILLER_97_28 ();
 FILLCELL_X2 FILLER_97_32 ();
 FILLCELL_X4 FILLER_97_41 ();
 FILLCELL_X2 FILLER_97_65 ();
 FILLCELL_X1 FILLER_97_67 ();
 FILLCELL_X1 FILLER_97_88 ();
 FILLCELL_X2 FILLER_97_110 ();
 FILLCELL_X1 FILLER_97_112 ();
 FILLCELL_X1 FILLER_97_132 ();
 FILLCELL_X4 FILLER_97_147 ();
 FILLCELL_X2 FILLER_97_151 ();
 FILLCELL_X1 FILLER_97_153 ();
 FILLCELL_X4 FILLER_97_181 ();
 FILLCELL_X2 FILLER_97_223 ();
 FILLCELL_X8 FILLER_97_245 ();
 FILLCELL_X4 FILLER_97_253 ();
 FILLCELL_X1 FILLER_97_257 ();
 FILLCELL_X8 FILLER_97_265 ();
 FILLCELL_X4 FILLER_97_273 ();
 FILLCELL_X8 FILLER_97_281 ();
 FILLCELL_X4 FILLER_97_292 ();
 FILLCELL_X8 FILLER_97_300 ();
 FILLCELL_X2 FILLER_97_311 ();
 FILLCELL_X1 FILLER_97_313 ();
 FILLCELL_X1 FILLER_97_318 ();
 FILLCELL_X4 FILLER_97_322 ();
 FILLCELL_X2 FILLER_97_326 ();
 FILLCELL_X4 FILLER_97_347 ();
 FILLCELL_X1 FILLER_97_351 ();
 FILLCELL_X4 FILLER_97_375 ();
 FILLCELL_X2 FILLER_97_379 ();
 FILLCELL_X4 FILLER_97_388 ();
 FILLCELL_X1 FILLER_97_392 ();
 FILLCELL_X2 FILLER_97_417 ();
 FILLCELL_X2 FILLER_97_427 ();
 FILLCELL_X2 FILLER_97_449 ();
 FILLCELL_X4 FILLER_97_465 ();
 FILLCELL_X2 FILLER_97_480 ();
 FILLCELL_X4 FILLER_97_489 ();
 FILLCELL_X4 FILLER_97_533 ();
 FILLCELL_X8 FILLER_97_540 ();
 FILLCELL_X2 FILLER_97_548 ();
 FILLCELL_X4 FILLER_97_570 ();
 FILLCELL_X2 FILLER_97_603 ();
 FILLCELL_X1 FILLER_97_632 ();
 FILLCELL_X2 FILLER_97_647 ();
 FILLCELL_X1 FILLER_97_649 ();
 FILLCELL_X2 FILLER_97_669 ();
 FILLCELL_X1 FILLER_97_678 ();
 FILLCELL_X1 FILLER_97_690 ();
 FILLCELL_X1 FILLER_97_698 ();
 FILLCELL_X4 FILLER_97_713 ();
 FILLCELL_X2 FILLER_97_717 ();
 FILLCELL_X1 FILLER_97_719 ();
 FILLCELL_X4 FILLER_97_738 ();
 FILLCELL_X1 FILLER_97_742 ();
 FILLCELL_X4 FILLER_97_747 ();
 FILLCELL_X2 FILLER_97_751 ();
 FILLCELL_X1 FILLER_97_753 ();
 FILLCELL_X2 FILLER_97_768 ();
 FILLCELL_X4 FILLER_97_781 ();
 FILLCELL_X1 FILLER_97_785 ();
 FILLCELL_X1 FILLER_97_796 ();
 FILLCELL_X8 FILLER_97_824 ();
 FILLCELL_X4 FILLER_97_837 ();
 FILLCELL_X2 FILLER_97_841 ();
 FILLCELL_X1 FILLER_97_843 ();
 FILLCELL_X2 FILLER_97_879 ();
 FILLCELL_X1 FILLER_97_881 ();
 FILLCELL_X1 FILLER_97_907 ();
 FILLCELL_X4 FILLER_97_921 ();
 FILLCELL_X2 FILLER_97_928 ();
 FILLCELL_X1 FILLER_97_939 ();
 FILLCELL_X1 FILLER_97_949 ();
 FILLCELL_X8 FILLER_97_954 ();
 FILLCELL_X2 FILLER_97_962 ();
 FILLCELL_X1 FILLER_97_964 ();
 FILLCELL_X8 FILLER_97_972 ();
 FILLCELL_X8 FILLER_97_987 ();
 FILLCELL_X4 FILLER_97_995 ();
 FILLCELL_X1 FILLER_97_999 ();
 FILLCELL_X4 FILLER_97_1007 ();
 FILLCELL_X1 FILLER_97_1011 ();
 FILLCELL_X2 FILLER_97_1041 ();
 FILLCELL_X1 FILLER_97_1043 ();
 FILLCELL_X16 FILLER_97_1071 ();
 FILLCELL_X1 FILLER_97_1087 ();
 FILLCELL_X8 FILLER_97_1127 ();
 FILLCELL_X2 FILLER_97_1135 ();
 FILLCELL_X1 FILLER_97_1137 ();
 FILLCELL_X4 FILLER_97_1172 ();
 FILLCELL_X4 FILLER_97_1212 ();
 FILLCELL_X1 FILLER_97_1216 ();
 FILLCELL_X2 FILLER_97_1221 ();
 FILLCELL_X1 FILLER_97_1223 ();
 FILLCELL_X2 FILLER_97_1250 ();
 FILLCELL_X1 FILLER_98_21 ();
 FILLCELL_X4 FILLER_98_43 ();
 FILLCELL_X2 FILLER_98_47 ();
 FILLCELL_X8 FILLER_98_56 ();
 FILLCELL_X2 FILLER_98_64 ();
 FILLCELL_X1 FILLER_98_66 ();
 FILLCELL_X8 FILLER_98_74 ();
 FILLCELL_X2 FILLER_98_82 ();
 FILLCELL_X1 FILLER_98_84 ();
 FILLCELL_X8 FILLER_98_92 ();
 FILLCELL_X4 FILLER_98_100 ();
 FILLCELL_X2 FILLER_98_104 ();
 FILLCELL_X1 FILLER_98_106 ();
 FILLCELL_X4 FILLER_98_127 ();
 FILLCELL_X4 FILLER_98_158 ();
 FILLCELL_X2 FILLER_98_162 ();
 FILLCELL_X2 FILLER_98_171 ();
 FILLCELL_X4 FILLER_98_176 ();
 FILLCELL_X8 FILLER_98_191 ();
 FILLCELL_X1 FILLER_98_199 ();
 FILLCELL_X2 FILLER_98_208 ();
 FILLCELL_X1 FILLER_98_210 ();
 FILLCELL_X1 FILLER_98_218 ();
 FILLCELL_X8 FILLER_98_226 ();
 FILLCELL_X2 FILLER_98_234 ();
 FILLCELL_X1 FILLER_98_243 ();
 FILLCELL_X1 FILLER_98_271 ();
 FILLCELL_X2 FILLER_98_292 ();
 FILLCELL_X1 FILLER_98_314 ();
 FILLCELL_X2 FILLER_98_320 ();
 FILLCELL_X16 FILLER_98_336 ();
 FILLCELL_X1 FILLER_98_352 ();
 FILLCELL_X8 FILLER_98_364 ();
 FILLCELL_X4 FILLER_98_372 ();
 FILLCELL_X2 FILLER_98_376 ();
 FILLCELL_X1 FILLER_98_378 ();
 FILLCELL_X4 FILLER_98_410 ();
 FILLCELL_X2 FILLER_98_414 ();
 FILLCELL_X1 FILLER_98_416 ();
 FILLCELL_X8 FILLER_98_420 ();
 FILLCELL_X4 FILLER_98_428 ();
 FILLCELL_X2 FILLER_98_432 ();
 FILLCELL_X1 FILLER_98_434 ();
 FILLCELL_X2 FILLER_98_446 ();
 FILLCELL_X2 FILLER_98_477 ();
 FILLCELL_X2 FILLER_98_486 ();
 FILLCELL_X2 FILLER_98_495 ();
 FILLCELL_X8 FILLER_98_500 ();
 FILLCELL_X2 FILLER_98_508 ();
 FILLCELL_X1 FILLER_98_510 ();
 FILLCELL_X8 FILLER_98_519 ();
 FILLCELL_X4 FILLER_98_554 ();
 FILLCELL_X16 FILLER_98_598 ();
 FILLCELL_X2 FILLER_98_614 ();
 FILLCELL_X1 FILLER_98_616 ();
 FILLCELL_X8 FILLER_98_632 ();
 FILLCELL_X2 FILLER_98_640 ();
 FILLCELL_X2 FILLER_98_651 ();
 FILLCELL_X1 FILLER_98_674 ();
 FILLCELL_X1 FILLER_98_684 ();
 FILLCELL_X2 FILLER_98_701 ();
 FILLCELL_X1 FILLER_98_703 ();
 FILLCELL_X16 FILLER_98_711 ();
 FILLCELL_X1 FILLER_98_727 ();
 FILLCELL_X2 FILLER_98_732 ();
 FILLCELL_X4 FILLER_98_738 ();
 FILLCELL_X1 FILLER_98_742 ();
 FILLCELL_X1 FILLER_98_768 ();
 FILLCELL_X4 FILLER_98_788 ();
 FILLCELL_X2 FILLER_98_811 ();
 FILLCELL_X4 FILLER_98_826 ();
 FILLCELL_X1 FILLER_98_830 ();
 FILLCELL_X2 FILLER_98_843 ();
 FILLCELL_X4 FILLER_98_874 ();
 FILLCELL_X2 FILLER_98_882 ();
 FILLCELL_X1 FILLER_98_884 ();
 FILLCELL_X2 FILLER_98_893 ();
 FILLCELL_X1 FILLER_98_899 ();
 FILLCELL_X2 FILLER_98_904 ();
 FILLCELL_X1 FILLER_98_906 ();
 FILLCELL_X8 FILLER_98_915 ();
 FILLCELL_X4 FILLER_98_923 ();
 FILLCELL_X1 FILLER_98_927 ();
 FILLCELL_X2 FILLER_98_931 ();
 FILLCELL_X4 FILLER_98_936 ();
 FILLCELL_X2 FILLER_98_940 ();
 FILLCELL_X2 FILLER_98_945 ();
 FILLCELL_X1 FILLER_98_947 ();
 FILLCELL_X4 FILLER_98_955 ();
 FILLCELL_X2 FILLER_98_959 ();
 FILLCELL_X4 FILLER_98_1025 ();
 FILLCELL_X2 FILLER_98_1029 ();
 FILLCELL_X8 FILLER_98_1049 ();
 FILLCELL_X4 FILLER_98_1057 ();
 FILLCELL_X1 FILLER_98_1061 ();
 FILLCELL_X16 FILLER_98_1069 ();
 FILLCELL_X8 FILLER_98_1085 ();
 FILLCELL_X2 FILLER_98_1093 ();
 FILLCELL_X2 FILLER_98_1100 ();
 FILLCELL_X4 FILLER_98_1115 ();
 FILLCELL_X16 FILLER_98_1160 ();
 FILLCELL_X8 FILLER_98_1176 ();
 FILLCELL_X4 FILLER_98_1184 ();
 FILLCELL_X2 FILLER_98_1188 ();
 FILLCELL_X1 FILLER_98_1190 ();
 FILLCELL_X4 FILLER_98_1198 ();
 FILLCELL_X2 FILLER_98_1202 ();
 FILLCELL_X1 FILLER_98_1222 ();
 FILLCELL_X8 FILLER_98_1229 ();
 FILLCELL_X2 FILLER_98_1237 ();
 FILLCELL_X8 FILLER_98_1246 ();
 FILLCELL_X1 FILLER_98_1254 ();
 FILLCELL_X8 FILLER_99_1 ();
 FILLCELL_X4 FILLER_99_9 ();
 FILLCELL_X8 FILLER_99_21 ();
 FILLCELL_X4 FILLER_99_29 ();
 FILLCELL_X1 FILLER_99_33 ();
 FILLCELL_X4 FILLER_99_61 ();
 FILLCELL_X8 FILLER_99_120 ();
 FILLCELL_X2 FILLER_99_128 ();
 FILLCELL_X8 FILLER_99_137 ();
 FILLCELL_X4 FILLER_99_145 ();
 FILLCELL_X1 FILLER_99_149 ();
 FILLCELL_X8 FILLER_99_157 ();
 FILLCELL_X2 FILLER_99_165 ();
 FILLCELL_X16 FILLER_99_187 ();
 FILLCELL_X4 FILLER_99_203 ();
 FILLCELL_X1 FILLER_99_207 ();
 FILLCELL_X8 FILLER_99_229 ();
 FILLCELL_X2 FILLER_99_237 ();
 FILLCELL_X2 FILLER_99_253 ();
 FILLCELL_X1 FILLER_99_255 ();
 FILLCELL_X2 FILLER_99_270 ();
 FILLCELL_X1 FILLER_99_272 ();
 FILLCELL_X1 FILLER_99_280 ();
 FILLCELL_X8 FILLER_99_288 ();
 FILLCELL_X4 FILLER_99_296 ();
 FILLCELL_X1 FILLER_99_300 ();
 FILLCELL_X2 FILLER_99_305 ();
 FILLCELL_X1 FILLER_99_307 ();
 FILLCELL_X2 FILLER_99_311 ();
 FILLCELL_X1 FILLER_99_313 ();
 FILLCELL_X4 FILLER_99_319 ();
 FILLCELL_X2 FILLER_99_323 ();
 FILLCELL_X4 FILLER_99_332 ();
 FILLCELL_X2 FILLER_99_336 ();
 FILLCELL_X4 FILLER_99_345 ();
 FILLCELL_X2 FILLER_99_369 ();
 FILLCELL_X2 FILLER_99_390 ();
 FILLCELL_X8 FILLER_99_410 ();
 FILLCELL_X4 FILLER_99_440 ();
 FILLCELL_X2 FILLER_99_444 ();
 FILLCELL_X2 FILLER_99_474 ();
 FILLCELL_X1 FILLER_99_505 ();
 FILLCELL_X1 FILLER_99_511 ();
 FILLCELL_X1 FILLER_99_516 ();
 FILLCELL_X8 FILLER_99_520 ();
 FILLCELL_X2 FILLER_99_528 ();
 FILLCELL_X1 FILLER_99_530 ();
 FILLCELL_X8 FILLER_99_558 ();
 FILLCELL_X4 FILLER_99_569 ();
 FILLCELL_X1 FILLER_99_573 ();
 FILLCELL_X8 FILLER_99_585 ();
 FILLCELL_X4 FILLER_99_593 ();
 FILLCELL_X2 FILLER_99_597 ();
 FILLCELL_X8 FILLER_99_620 ();
 FILLCELL_X2 FILLER_99_628 ();
 FILLCELL_X16 FILLER_99_640 ();
 FILLCELL_X8 FILLER_99_656 ();
 FILLCELL_X1 FILLER_99_664 ();
 FILLCELL_X16 FILLER_99_679 ();
 FILLCELL_X1 FILLER_99_695 ();
 FILLCELL_X2 FILLER_99_728 ();
 FILLCELL_X1 FILLER_99_730 ();
 FILLCELL_X2 FILLER_99_738 ();
 FILLCELL_X1 FILLER_99_740 ();
 FILLCELL_X1 FILLER_99_745 ();
 FILLCELL_X4 FILLER_99_754 ();
 FILLCELL_X1 FILLER_99_758 ();
 FILLCELL_X2 FILLER_99_775 ();
 FILLCELL_X2 FILLER_99_791 ();
 FILLCELL_X4 FILLER_99_796 ();
 FILLCELL_X1 FILLER_99_800 ();
 FILLCELL_X4 FILLER_99_807 ();
 FILLCELL_X2 FILLER_99_811 ();
 FILLCELL_X1 FILLER_99_813 ();
 FILLCELL_X1 FILLER_99_820 ();
 FILLCELL_X1 FILLER_99_832 ();
 FILLCELL_X16 FILLER_99_853 ();
 FILLCELL_X4 FILLER_99_869 ();
 FILLCELL_X2 FILLER_99_873 ();
 FILLCELL_X1 FILLER_99_875 ();
 FILLCELL_X1 FILLER_99_892 ();
 FILLCELL_X1 FILLER_99_897 ();
 FILLCELL_X1 FILLER_99_908 ();
 FILLCELL_X1 FILLER_99_913 ();
 FILLCELL_X2 FILLER_99_921 ();
 FILLCELL_X2 FILLER_99_926 ();
 FILLCELL_X8 FILLER_99_931 ();
 FILLCELL_X4 FILLER_99_939 ();
 FILLCELL_X2 FILLER_99_943 ();
 FILLCELL_X1 FILLER_99_945 ();
 FILLCELL_X16 FILLER_99_964 ();
 FILLCELL_X8 FILLER_99_980 ();
 FILLCELL_X4 FILLER_99_988 ();
 FILLCELL_X2 FILLER_99_992 ();
 FILLCELL_X8 FILLER_99_998 ();
 FILLCELL_X1 FILLER_99_1006 ();
 FILLCELL_X4 FILLER_99_1024 ();
 FILLCELL_X2 FILLER_99_1028 ();
 FILLCELL_X1 FILLER_99_1030 ();
 FILLCELL_X16 FILLER_99_1045 ();
 FILLCELL_X8 FILLER_99_1061 ();
 FILLCELL_X2 FILLER_99_1069 ();
 FILLCELL_X1 FILLER_99_1071 ();
 FILLCELL_X8 FILLER_99_1075 ();
 FILLCELL_X2 FILLER_99_1083 ();
 FILLCELL_X1 FILLER_99_1085 ();
 FILLCELL_X8 FILLER_99_1093 ();
 FILLCELL_X1 FILLER_99_1101 ();
 FILLCELL_X2 FILLER_99_1105 ();
 FILLCELL_X8 FILLER_99_1110 ();
 FILLCELL_X2 FILLER_99_1118 ();
 FILLCELL_X1 FILLER_99_1120 ();
 FILLCELL_X8 FILLER_99_1126 ();
 FILLCELL_X1 FILLER_99_1134 ();
 FILLCELL_X4 FILLER_99_1141 ();
 FILLCELL_X1 FILLER_99_1145 ();
 FILLCELL_X4 FILLER_99_1149 ();
 FILLCELL_X1 FILLER_99_1162 ();
 FILLCELL_X2 FILLER_99_1170 ();
 FILLCELL_X1 FILLER_99_1172 ();
 FILLCELL_X2 FILLER_99_1189 ();
 FILLCELL_X1 FILLER_99_1191 ();
 FILLCELL_X1 FILLER_99_1205 ();
 FILLCELL_X8 FILLER_99_1230 ();
 FILLCELL_X1 FILLER_99_1238 ();
 FILLCELL_X2 FILLER_99_1249 ();
 FILLCELL_X1 FILLER_99_1254 ();
 FILLCELL_X4 FILLER_100_1 ();
 FILLCELL_X8 FILLER_100_32 ();
 FILLCELL_X1 FILLER_100_40 ();
 FILLCELL_X16 FILLER_100_48 ();
 FILLCELL_X4 FILLER_100_64 ();
 FILLCELL_X2 FILLER_100_68 ();
 FILLCELL_X1 FILLER_100_84 ();
 FILLCELL_X1 FILLER_100_92 ();
 FILLCELL_X2 FILLER_100_100 ();
 FILLCELL_X2 FILLER_100_156 ();
 FILLCELL_X4 FILLER_100_165 ();
 FILLCELL_X2 FILLER_100_169 ();
 FILLCELL_X1 FILLER_100_171 ();
 FILLCELL_X2 FILLER_100_185 ();
 FILLCELL_X1 FILLER_100_187 ();
 FILLCELL_X1 FILLER_100_202 ();
 FILLCELL_X4 FILLER_100_210 ();
 FILLCELL_X2 FILLER_100_214 ();
 FILLCELL_X1 FILLER_100_216 ();
 FILLCELL_X8 FILLER_100_224 ();
 FILLCELL_X1 FILLER_100_232 ();
 FILLCELL_X2 FILLER_100_254 ();
 FILLCELL_X1 FILLER_100_256 ();
 FILLCELL_X8 FILLER_100_283 ();
 FILLCELL_X4 FILLER_100_291 ();
 FILLCELL_X2 FILLER_100_295 ();
 FILLCELL_X4 FILLER_100_317 ();
 FILLCELL_X4 FILLER_100_348 ();
 FILLCELL_X2 FILLER_100_352 ();
 FILLCELL_X4 FILLER_100_361 ();
 FILLCELL_X4 FILLER_100_388 ();
 FILLCELL_X8 FILLER_100_399 ();
 FILLCELL_X4 FILLER_100_407 ();
 FILLCELL_X2 FILLER_100_411 ();
 FILLCELL_X1 FILLER_100_413 ();
 FILLCELL_X4 FILLER_100_421 ();
 FILLCELL_X1 FILLER_100_436 ();
 FILLCELL_X2 FILLER_100_444 ();
 FILLCELL_X1 FILLER_100_446 ();
 FILLCELL_X8 FILLER_100_450 ();
 FILLCELL_X8 FILLER_100_474 ();
 FILLCELL_X1 FILLER_100_482 ();
 FILLCELL_X8 FILLER_100_490 ();
 FILLCELL_X4 FILLER_100_498 ();
 FILLCELL_X2 FILLER_100_502 ();
 FILLCELL_X1 FILLER_100_504 ();
 FILLCELL_X4 FILLER_100_541 ();
 FILLCELL_X1 FILLER_100_545 ();
 FILLCELL_X8 FILLER_100_587 ();
 FILLCELL_X8 FILLER_100_612 ();
 FILLCELL_X4 FILLER_100_620 ();
 FILLCELL_X2 FILLER_100_635 ();
 FILLCELL_X1 FILLER_100_637 ();
 FILLCELL_X2 FILLER_100_642 ();
 FILLCELL_X1 FILLER_100_644 ();
 FILLCELL_X4 FILLER_100_654 ();
 FILLCELL_X2 FILLER_100_658 ();
 FILLCELL_X1 FILLER_100_660 ();
 FILLCELL_X2 FILLER_100_674 ();
 FILLCELL_X1 FILLER_100_680 ();
 FILLCELL_X32 FILLER_100_686 ();
 FILLCELL_X8 FILLER_100_718 ();
 FILLCELL_X4 FILLER_100_731 ();
 FILLCELL_X1 FILLER_100_735 ();
 FILLCELL_X2 FILLER_100_741 ();
 FILLCELL_X1 FILLER_100_743 ();
 FILLCELL_X2 FILLER_100_749 ();
 FILLCELL_X2 FILLER_100_763 ();
 FILLCELL_X1 FILLER_100_765 ();
 FILLCELL_X2 FILLER_100_791 ();
 FILLCELL_X1 FILLER_100_793 ();
 FILLCELL_X1 FILLER_100_801 ();
 FILLCELL_X1 FILLER_100_809 ();
 FILLCELL_X2 FILLER_100_818 ();
 FILLCELL_X8 FILLER_100_839 ();
 FILLCELL_X4 FILLER_100_847 ();
 FILLCELL_X4 FILLER_100_884 ();
 FILLCELL_X1 FILLER_100_888 ();
 FILLCELL_X1 FILLER_100_896 ();
 FILLCELL_X1 FILLER_100_906 ();
 FILLCELL_X1 FILLER_100_924 ();
 FILLCELL_X8 FILLER_100_936 ();
 FILLCELL_X4 FILLER_100_944 ();
 FILLCELL_X2 FILLER_100_948 ();
 FILLCELL_X16 FILLER_100_963 ();
 FILLCELL_X1 FILLER_100_986 ();
 FILLCELL_X1 FILLER_100_996 ();
 FILLCELL_X2 FILLER_100_1004 ();
 FILLCELL_X1 FILLER_100_1015 ();
 FILLCELL_X4 FILLER_100_1031 ();
 FILLCELL_X1 FILLER_100_1035 ();
 FILLCELL_X8 FILLER_100_1049 ();
 FILLCELL_X2 FILLER_100_1077 ();
 FILLCELL_X1 FILLER_100_1102 ();
 FILLCELL_X4 FILLER_100_1110 ();
 FILLCELL_X1 FILLER_100_1114 ();
 FILLCELL_X1 FILLER_100_1147 ();
 FILLCELL_X1 FILLER_100_1154 ();
 FILLCELL_X2 FILLER_100_1160 ();
 FILLCELL_X4 FILLER_100_1166 ();
 FILLCELL_X1 FILLER_100_1170 ();
 FILLCELL_X4 FILLER_100_1209 ();
 FILLCELL_X1 FILLER_100_1216 ();
 FILLCELL_X2 FILLER_100_1221 ();
 FILLCELL_X2 FILLER_100_1228 ();
 FILLCELL_X2 FILLER_100_1233 ();
 FILLCELL_X2 FILLER_100_1252 ();
 FILLCELL_X1 FILLER_100_1254 ();
 FILLCELL_X4 FILLER_101_1 ();
 FILLCELL_X1 FILLER_101_5 ();
 FILLCELL_X16 FILLER_101_47 ();
 FILLCELL_X8 FILLER_101_63 ();
 FILLCELL_X32 FILLER_101_106 ();
 FILLCELL_X8 FILLER_101_138 ();
 FILLCELL_X2 FILLER_101_160 ();
 FILLCELL_X8 FILLER_101_191 ();
 FILLCELL_X2 FILLER_101_206 ();
 FILLCELL_X8 FILLER_101_228 ();
 FILLCELL_X2 FILLER_101_236 ();
 FILLCELL_X1 FILLER_101_238 ();
 FILLCELL_X2 FILLER_101_243 ();
 FILLCELL_X1 FILLER_101_245 ();
 FILLCELL_X8 FILLER_101_249 ();
 FILLCELL_X1 FILLER_101_262 ();
 FILLCELL_X8 FILLER_101_266 ();
 FILLCELL_X4 FILLER_101_279 ();
 FILLCELL_X8 FILLER_101_303 ();
 FILLCELL_X1 FILLER_101_325 ();
 FILLCELL_X2 FILLER_101_333 ();
 FILLCELL_X16 FILLER_101_342 ();
 FILLCELL_X1 FILLER_101_358 ();
 FILLCELL_X4 FILLER_101_373 ();
 FILLCELL_X2 FILLER_101_377 ();
 FILLCELL_X1 FILLER_101_379 ();
 FILLCELL_X1 FILLER_101_407 ();
 FILLCELL_X8 FILLER_101_448 ();
 FILLCELL_X4 FILLER_101_456 ();
 FILLCELL_X2 FILLER_101_460 ();
 FILLCELL_X8 FILLER_101_489 ();
 FILLCELL_X4 FILLER_101_497 ();
 FILLCELL_X1 FILLER_101_501 ();
 FILLCELL_X2 FILLER_101_515 ();
 FILLCELL_X4 FILLER_101_545 ();
 FILLCELL_X8 FILLER_101_563 ();
 FILLCELL_X4 FILLER_101_571 ();
 FILLCELL_X1 FILLER_101_575 ();
 FILLCELL_X2 FILLER_101_579 ();
 FILLCELL_X2 FILLER_101_608 ();
 FILLCELL_X4 FILLER_101_617 ();
 FILLCELL_X4 FILLER_101_642 ();
 FILLCELL_X2 FILLER_101_651 ();
 FILLCELL_X1 FILLER_101_653 ();
 FILLCELL_X4 FILLER_101_678 ();
 FILLCELL_X1 FILLER_101_682 ();
 FILLCELL_X4 FILLER_101_695 ();
 FILLCELL_X1 FILLER_101_699 ();
 FILLCELL_X4 FILLER_101_704 ();
 FILLCELL_X2 FILLER_101_708 ();
 FILLCELL_X4 FILLER_101_721 ();
 FILLCELL_X2 FILLER_101_725 ();
 FILLCELL_X8 FILLER_101_738 ();
 FILLCELL_X2 FILLER_101_746 ();
 FILLCELL_X1 FILLER_101_748 ();
 FILLCELL_X4 FILLER_101_757 ();
 FILLCELL_X1 FILLER_101_761 ();
 FILLCELL_X2 FILLER_101_771 ();
 FILLCELL_X4 FILLER_101_775 ();
 FILLCELL_X2 FILLER_101_779 ();
 FILLCELL_X1 FILLER_101_781 ();
 FILLCELL_X1 FILLER_101_804 ();
 FILLCELL_X4 FILLER_101_817 ();
 FILLCELL_X2 FILLER_101_821 ();
 FILLCELL_X1 FILLER_101_823 ();
 FILLCELL_X4 FILLER_101_841 ();
 FILLCELL_X8 FILLER_101_854 ();
 FILLCELL_X4 FILLER_101_862 ();
 FILLCELL_X1 FILLER_101_866 ();
 FILLCELL_X4 FILLER_101_870 ();
 FILLCELL_X1 FILLER_101_891 ();
 FILLCELL_X8 FILLER_101_895 ();
 FILLCELL_X2 FILLER_101_903 ();
 FILLCELL_X1 FILLER_101_905 ();
 FILLCELL_X1 FILLER_101_913 ();
 FILLCELL_X4 FILLER_101_924 ();
 FILLCELL_X1 FILLER_101_928 ();
 FILLCELL_X8 FILLER_101_936 ();
 FILLCELL_X4 FILLER_101_944 ();
 FILLCELL_X2 FILLER_101_948 ();
 FILLCELL_X1 FILLER_101_950 ();
 FILLCELL_X1 FILLER_101_960 ();
 FILLCELL_X1 FILLER_101_971 ();
 FILLCELL_X1 FILLER_101_976 ();
 FILLCELL_X1 FILLER_101_981 ();
 FILLCELL_X32 FILLER_101_997 ();
 FILLCELL_X2 FILLER_101_1029 ();
 FILLCELL_X16 FILLER_101_1037 ();
 FILLCELL_X8 FILLER_101_1053 ();
 FILLCELL_X2 FILLER_101_1082 ();
 FILLCELL_X1 FILLER_101_1084 ();
 FILLCELL_X16 FILLER_101_1088 ();
 FILLCELL_X4 FILLER_101_1119 ();
 FILLCELL_X2 FILLER_101_1123 ();
 FILLCELL_X1 FILLER_101_1125 ();
 FILLCELL_X8 FILLER_101_1165 ();
 FILLCELL_X2 FILLER_101_1173 ();
 FILLCELL_X1 FILLER_101_1175 ();
 FILLCELL_X4 FILLER_101_1183 ();
 FILLCELL_X8 FILLER_101_1192 ();
 FILLCELL_X2 FILLER_101_1248 ();
 FILLCELL_X2 FILLER_101_1253 ();
 FILLCELL_X4 FILLER_102_1 ();
 FILLCELL_X1 FILLER_102_5 ();
 FILLCELL_X8 FILLER_102_13 ();
 FILLCELL_X4 FILLER_102_21 ();
 FILLCELL_X1 FILLER_102_25 ();
 FILLCELL_X2 FILLER_102_33 ();
 FILLCELL_X2 FILLER_102_42 ();
 FILLCELL_X1 FILLER_102_44 ();
 FILLCELL_X4 FILLER_102_65 ();
 FILLCELL_X1 FILLER_102_69 ();
 FILLCELL_X4 FILLER_102_77 ();
 FILLCELL_X1 FILLER_102_81 ();
 FILLCELL_X4 FILLER_102_89 ();
 FILLCELL_X2 FILLER_102_107 ();
 FILLCELL_X8 FILLER_102_143 ();
 FILLCELL_X4 FILLER_102_151 ();
 FILLCELL_X2 FILLER_102_155 ();
 FILLCELL_X4 FILLER_102_183 ();
 FILLCELL_X1 FILLER_102_187 ();
 FILLCELL_X1 FILLER_102_208 ();
 FILLCELL_X8 FILLER_102_223 ();
 FILLCELL_X1 FILLER_102_231 ();
 FILLCELL_X2 FILLER_102_299 ();
 FILLCELL_X2 FILLER_102_321 ();
 FILLCELL_X1 FILLER_102_323 ();
 FILLCELL_X16 FILLER_102_331 ();
 FILLCELL_X2 FILLER_102_347 ();
 FILLCELL_X4 FILLER_102_396 ();
 FILLCELL_X2 FILLER_102_400 ();
 FILLCELL_X1 FILLER_102_402 ();
 FILLCELL_X4 FILLER_102_410 ();
 FILLCELL_X4 FILLER_102_421 ();
 FILLCELL_X1 FILLER_102_425 ();
 FILLCELL_X8 FILLER_102_467 ();
 FILLCELL_X4 FILLER_102_475 ();
 FILLCELL_X2 FILLER_102_479 ();
 FILLCELL_X1 FILLER_102_481 ();
 FILLCELL_X4 FILLER_102_509 ();
 FILLCELL_X2 FILLER_102_513 ();
 FILLCELL_X1 FILLER_102_535 ();
 FILLCELL_X8 FILLER_102_543 ();
 FILLCELL_X1 FILLER_102_551 ();
 FILLCELL_X8 FILLER_102_579 ();
 FILLCELL_X2 FILLER_102_594 ();
 FILLCELL_X1 FILLER_102_596 ();
 FILLCELL_X2 FILLER_102_632 ();
 FILLCELL_X8 FILLER_102_641 ();
 FILLCELL_X4 FILLER_102_649 ();
 FILLCELL_X1 FILLER_102_684 ();
 FILLCELL_X4 FILLER_102_736 ();
 FILLCELL_X2 FILLER_102_740 ();
 FILLCELL_X1 FILLER_102_746 ();
 FILLCELL_X2 FILLER_102_751 ();
 FILLCELL_X4 FILLER_102_757 ();
 FILLCELL_X2 FILLER_102_765 ();
 FILLCELL_X16 FILLER_102_777 ();
 FILLCELL_X4 FILLER_102_793 ();
 FILLCELL_X2 FILLER_102_797 ();
 FILLCELL_X4 FILLER_102_810 ();
 FILLCELL_X1 FILLER_102_814 ();
 FILLCELL_X4 FILLER_102_820 ();
 FILLCELL_X8 FILLER_102_834 ();
 FILLCELL_X2 FILLER_102_842 ();
 FILLCELL_X1 FILLER_102_844 ();
 FILLCELL_X2 FILLER_102_855 ();
 FILLCELL_X1 FILLER_102_857 ();
 FILLCELL_X2 FILLER_102_860 ();
 FILLCELL_X4 FILLER_102_873 ();
 FILLCELL_X2 FILLER_102_895 ();
 FILLCELL_X8 FILLER_102_906 ();
 FILLCELL_X2 FILLER_102_914 ();
 FILLCELL_X4 FILLER_102_925 ();
 FILLCELL_X2 FILLER_102_929 ();
 FILLCELL_X1 FILLER_102_931 ();
 FILLCELL_X1 FILLER_102_983 ();
 FILLCELL_X1 FILLER_102_989 ();
 FILLCELL_X4 FILLER_102_1025 ();
 FILLCELL_X2 FILLER_102_1029 ();
 FILLCELL_X2 FILLER_102_1042 ();
 FILLCELL_X1 FILLER_102_1044 ();
 FILLCELL_X8 FILLER_102_1052 ();
 FILLCELL_X2 FILLER_102_1060 ();
 FILLCELL_X1 FILLER_102_1062 ();
 FILLCELL_X2 FILLER_102_1076 ();
 FILLCELL_X4 FILLER_102_1084 ();
 FILLCELL_X2 FILLER_102_1088 ();
 FILLCELL_X8 FILLER_102_1116 ();
 FILLCELL_X4 FILLER_102_1124 ();
 FILLCELL_X4 FILLER_102_1139 ();
 FILLCELL_X2 FILLER_102_1143 ();
 FILLCELL_X1 FILLER_102_1145 ();
 FILLCELL_X2 FILLER_102_1172 ();
 FILLCELL_X1 FILLER_102_1194 ();
 FILLCELL_X16 FILLER_102_1202 ();
 FILLCELL_X1 FILLER_102_1218 ();
 FILLCELL_X8 FILLER_102_1226 ();
 FILLCELL_X4 FILLER_102_1234 ();
 FILLCELL_X4 FILLER_102_1248 ();
 FILLCELL_X8 FILLER_103_35 ();
 FILLCELL_X4 FILLER_103_43 ();
 FILLCELL_X2 FILLER_103_47 ();
 FILLCELL_X1 FILLER_103_49 ();
 FILLCELL_X1 FILLER_103_77 ();
 FILLCELL_X2 FILLER_103_92 ();
 FILLCELL_X1 FILLER_103_94 ();
 FILLCELL_X4 FILLER_103_109 ();
 FILLCELL_X2 FILLER_103_113 ();
 FILLCELL_X1 FILLER_103_115 ();
 FILLCELL_X8 FILLER_103_123 ();
 FILLCELL_X4 FILLER_103_131 ();
 FILLCELL_X4 FILLER_103_183 ();
 FILLCELL_X1 FILLER_103_187 ();
 FILLCELL_X1 FILLER_103_211 ();
 FILLCELL_X2 FILLER_103_219 ();
 FILLCELL_X2 FILLER_103_228 ();
 FILLCELL_X8 FILLER_103_237 ();
 FILLCELL_X2 FILLER_103_245 ();
 FILLCELL_X1 FILLER_103_247 ();
 FILLCELL_X4 FILLER_103_251 ();
 FILLCELL_X2 FILLER_103_255 ();
 FILLCELL_X4 FILLER_103_261 ();
 FILLCELL_X4 FILLER_103_286 ();
 FILLCELL_X2 FILLER_103_290 ();
 FILLCELL_X1 FILLER_103_292 ();
 FILLCELL_X2 FILLER_103_297 ();
 FILLCELL_X1 FILLER_103_299 ();
 FILLCELL_X8 FILLER_103_303 ();
 FILLCELL_X4 FILLER_103_311 ();
 FILLCELL_X2 FILLER_103_315 ();
 FILLCELL_X1 FILLER_103_317 ();
 FILLCELL_X1 FILLER_103_332 ();
 FILLCELL_X1 FILLER_103_351 ();
 FILLCELL_X4 FILLER_103_359 ();
 FILLCELL_X2 FILLER_103_363 ();
 FILLCELL_X4 FILLER_103_385 ();
 FILLCELL_X1 FILLER_103_389 ();
 FILLCELL_X1 FILLER_103_410 ();
 FILLCELL_X8 FILLER_103_438 ();
 FILLCELL_X4 FILLER_103_453 ();
 FILLCELL_X2 FILLER_103_457 ();
 FILLCELL_X4 FILLER_103_473 ();
 FILLCELL_X2 FILLER_103_477 ();
 FILLCELL_X8 FILLER_103_483 ();
 FILLCELL_X2 FILLER_103_491 ();
 FILLCELL_X4 FILLER_103_504 ();
 FILLCELL_X4 FILLER_103_535 ();
 FILLCELL_X1 FILLER_103_539 ();
 FILLCELL_X4 FILLER_103_554 ();
 FILLCELL_X2 FILLER_103_558 ();
 FILLCELL_X1 FILLER_103_560 ();
 FILLCELL_X8 FILLER_103_566 ();
 FILLCELL_X2 FILLER_103_574 ();
 FILLCELL_X1 FILLER_103_576 ();
 FILLCELL_X8 FILLER_103_638 ();
 FILLCELL_X4 FILLER_103_646 ();
 FILLCELL_X8 FILLER_103_663 ();
 FILLCELL_X2 FILLER_103_671 ();
 FILLCELL_X1 FILLER_103_673 ();
 FILLCELL_X4 FILLER_103_705 ();
 FILLCELL_X1 FILLER_103_709 ();
 FILLCELL_X4 FILLER_103_713 ();
 FILLCELL_X1 FILLER_103_717 ();
 FILLCELL_X4 FILLER_103_727 ();
 FILLCELL_X2 FILLER_103_731 ();
 FILLCELL_X1 FILLER_103_733 ();
 FILLCELL_X4 FILLER_103_738 ();
 FILLCELL_X8 FILLER_103_757 ();
 FILLCELL_X1 FILLER_103_765 ();
 FILLCELL_X4 FILLER_103_772 ();
 FILLCELL_X1 FILLER_103_776 ();
 FILLCELL_X1 FILLER_103_817 ();
 FILLCELL_X4 FILLER_103_824 ();
 FILLCELL_X1 FILLER_103_828 ();
 FILLCELL_X4 FILLER_103_837 ();
 FILLCELL_X8 FILLER_103_859 ();
 FILLCELL_X1 FILLER_103_867 ();
 FILLCELL_X2 FILLER_103_894 ();
 FILLCELL_X1 FILLER_103_940 ();
 FILLCELL_X2 FILLER_103_946 ();
 FILLCELL_X1 FILLER_103_955 ();
 FILLCELL_X2 FILLER_103_961 ();
 FILLCELL_X1 FILLER_103_963 ();
 FILLCELL_X1 FILLER_103_968 ();
 FILLCELL_X1 FILLER_103_974 ();
 FILLCELL_X1 FILLER_103_988 ();
 FILLCELL_X2 FILLER_103_1005 ();
 FILLCELL_X1 FILLER_103_1007 ();
 FILLCELL_X1 FILLER_103_1020 ();
 FILLCELL_X1 FILLER_103_1031 ();
 FILLCELL_X1 FILLER_103_1036 ();
 FILLCELL_X1 FILLER_103_1044 ();
 FILLCELL_X4 FILLER_103_1051 ();
 FILLCELL_X4 FILLER_103_1070 ();
 FILLCELL_X1 FILLER_103_1074 ();
 FILLCELL_X4 FILLER_103_1099 ();
 FILLCELL_X1 FILLER_103_1112 ();
 FILLCELL_X2 FILLER_103_1138 ();
 FILLCELL_X1 FILLER_103_1140 ();
 FILLCELL_X2 FILLER_103_1192 ();
 FILLCELL_X1 FILLER_103_1194 ();
 FILLCELL_X2 FILLER_103_1231 ();
 FILLCELL_X1 FILLER_103_1233 ();
 FILLCELL_X1 FILLER_103_1241 ();
 FILLCELL_X2 FILLER_103_1252 ();
 FILLCELL_X1 FILLER_103_1254 ();
 FILLCELL_X4 FILLER_104_1 ();
 FILLCELL_X1 FILLER_104_5 ();
 FILLCELL_X8 FILLER_104_13 ();
 FILLCELL_X2 FILLER_104_48 ();
 FILLCELL_X1 FILLER_104_50 ();
 FILLCELL_X8 FILLER_104_99 ();
 FILLCELL_X4 FILLER_104_107 ();
 FILLCELL_X2 FILLER_104_111 ();
 FILLCELL_X1 FILLER_104_113 ();
 FILLCELL_X8 FILLER_104_141 ();
 FILLCELL_X4 FILLER_104_149 ();
 FILLCELL_X2 FILLER_104_153 ();
 FILLCELL_X1 FILLER_104_155 ();
 FILLCELL_X1 FILLER_104_170 ();
 FILLCELL_X2 FILLER_104_181 ();
 FILLCELL_X1 FILLER_104_186 ();
 FILLCELL_X2 FILLER_104_196 ();
 FILLCELL_X1 FILLER_104_198 ();
 FILLCELL_X1 FILLER_104_203 ();
 FILLCELL_X1 FILLER_104_229 ();
 FILLCELL_X1 FILLER_104_250 ();
 FILLCELL_X2 FILLER_104_285 ();
 FILLCELL_X1 FILLER_104_287 ();
 FILLCELL_X2 FILLER_104_308 ();
 FILLCELL_X2 FILLER_104_314 ();
 FILLCELL_X1 FILLER_104_316 ();
 FILLCELL_X2 FILLER_104_334 ();
 FILLCELL_X2 FILLER_104_343 ();
 FILLCELL_X4 FILLER_104_365 ();
 FILLCELL_X2 FILLER_104_369 ();
 FILLCELL_X1 FILLER_104_378 ();
 FILLCELL_X4 FILLER_104_400 ();
 FILLCELL_X2 FILLER_104_404 ();
 FILLCELL_X8 FILLER_104_411 ();
 FILLCELL_X4 FILLER_104_419 ();
 FILLCELL_X4 FILLER_104_437 ();
 FILLCELL_X2 FILLER_104_499 ();
 FILLCELL_X8 FILLER_104_513 ();
 FILLCELL_X2 FILLER_104_521 ();
 FILLCELL_X2 FILLER_104_550 ();
 FILLCELL_X1 FILLER_104_552 ();
 FILLCELL_X2 FILLER_104_580 ();
 FILLCELL_X16 FILLER_104_589 ();
 FILLCELL_X8 FILLER_104_605 ();
 FILLCELL_X4 FILLER_104_613 ();
 FILLCELL_X2 FILLER_104_617 ();
 FILLCELL_X1 FILLER_104_619 ();
 FILLCELL_X4 FILLER_104_627 ();
 FILLCELL_X16 FILLER_104_632 ();
 FILLCELL_X8 FILLER_104_648 ();
 FILLCELL_X4 FILLER_104_669 ();
 FILLCELL_X1 FILLER_104_673 ();
 FILLCELL_X1 FILLER_104_699 ();
 FILLCELL_X1 FILLER_104_704 ();
 FILLCELL_X1 FILLER_104_710 ();
 FILLCELL_X2 FILLER_104_716 ();
 FILLCELL_X2 FILLER_104_731 ();
 FILLCELL_X4 FILLER_104_737 ();
 FILLCELL_X2 FILLER_104_741 ();
 FILLCELL_X1 FILLER_104_743 ();
 FILLCELL_X1 FILLER_104_754 ();
 FILLCELL_X1 FILLER_104_765 ();
 FILLCELL_X1 FILLER_104_777 ();
 FILLCELL_X2 FILLER_104_804 ();
 FILLCELL_X1 FILLER_104_813 ();
 FILLCELL_X8 FILLER_104_855 ();
 FILLCELL_X4 FILLER_104_863 ();
 FILLCELL_X8 FILLER_104_871 ();
 FILLCELL_X1 FILLER_104_879 ();
 FILLCELL_X1 FILLER_104_897 ();
 FILLCELL_X2 FILLER_104_905 ();
 FILLCELL_X2 FILLER_104_920 ();
 FILLCELL_X1 FILLER_104_926 ();
 FILLCELL_X4 FILLER_104_980 ();
 FILLCELL_X1 FILLER_104_984 ();
 FILLCELL_X4 FILLER_104_988 ();
 FILLCELL_X2 FILLER_104_994 ();
 FILLCELL_X4 FILLER_104_998 ();
 FILLCELL_X1 FILLER_104_1023 ();
 FILLCELL_X2 FILLER_104_1026 ();
 FILLCELL_X1 FILLER_104_1035 ();
 FILLCELL_X8 FILLER_104_1042 ();
 FILLCELL_X2 FILLER_104_1055 ();
 FILLCELL_X1 FILLER_104_1057 ();
 FILLCELL_X2 FILLER_104_1068 ();
 FILLCELL_X1 FILLER_104_1070 ();
 FILLCELL_X16 FILLER_104_1090 ();
 FILLCELL_X1 FILLER_104_1106 ();
 FILLCELL_X2 FILLER_104_1118 ();
 FILLCELL_X1 FILLER_104_1120 ();
 FILLCELL_X4 FILLER_104_1123 ();
 FILLCELL_X1 FILLER_104_1127 ();
 FILLCELL_X1 FILLER_104_1134 ();
 FILLCELL_X1 FILLER_104_1139 ();
 FILLCELL_X1 FILLER_104_1154 ();
 FILLCELL_X2 FILLER_104_1166 ();
 FILLCELL_X1 FILLER_104_1168 ();
 FILLCELL_X4 FILLER_104_1177 ();
 FILLCELL_X1 FILLER_104_1210 ();
 FILLCELL_X1 FILLER_104_1215 ();
 FILLCELL_X2 FILLER_104_1253 ();
 FILLCELL_X8 FILLER_105_1 ();
 FILLCELL_X8 FILLER_105_41 ();
 FILLCELL_X4 FILLER_105_56 ();
 FILLCELL_X2 FILLER_105_60 ();
 FILLCELL_X4 FILLER_105_69 ();
 FILLCELL_X1 FILLER_105_114 ();
 FILLCELL_X2 FILLER_105_122 ();
 FILLCELL_X1 FILLER_105_124 ();
 FILLCELL_X4 FILLER_105_140 ();
 FILLCELL_X2 FILLER_105_144 ();
 FILLCELL_X1 FILLER_105_146 ();
 FILLCELL_X4 FILLER_105_157 ();
 FILLCELL_X2 FILLER_105_175 ();
 FILLCELL_X1 FILLER_105_177 ();
 FILLCELL_X2 FILLER_105_183 ();
 FILLCELL_X4 FILLER_105_192 ();
 FILLCELL_X1 FILLER_105_196 ();
 FILLCELL_X16 FILLER_105_220 ();
 FILLCELL_X4 FILLER_105_236 ();
 FILLCELL_X1 FILLER_105_244 ();
 FILLCELL_X8 FILLER_105_248 ();
 FILLCELL_X4 FILLER_105_260 ();
 FILLCELL_X4 FILLER_105_274 ();
 FILLCELL_X2 FILLER_105_278 ();
 FILLCELL_X1 FILLER_105_280 ();
 FILLCELL_X4 FILLER_105_291 ();
 FILLCELL_X2 FILLER_105_299 ();
 FILLCELL_X4 FILLER_105_331 ();
 FILLCELL_X2 FILLER_105_335 ();
 FILLCELL_X4 FILLER_105_343 ();
 FILLCELL_X2 FILLER_105_347 ();
 FILLCELL_X1 FILLER_105_349 ();
 FILLCELL_X4 FILLER_105_357 ();
 FILLCELL_X1 FILLER_105_361 ();
 FILLCELL_X16 FILLER_105_369 ();
 FILLCELL_X4 FILLER_105_385 ();
 FILLCELL_X1 FILLER_105_389 ();
 FILLCELL_X4 FILLER_105_397 ();
 FILLCELL_X2 FILLER_105_401 ();
 FILLCELL_X8 FILLER_105_417 ();
 FILLCELL_X1 FILLER_105_425 ();
 FILLCELL_X16 FILLER_105_433 ();
 FILLCELL_X8 FILLER_105_449 ();
 FILLCELL_X2 FILLER_105_457 ();
 FILLCELL_X1 FILLER_105_459 ();
 FILLCELL_X1 FILLER_105_467 ();
 FILLCELL_X8 FILLER_105_475 ();
 FILLCELL_X4 FILLER_105_483 ();
 FILLCELL_X1 FILLER_105_487 ();
 FILLCELL_X8 FILLER_105_491 ();
 FILLCELL_X2 FILLER_105_499 ();
 FILLCELL_X1 FILLER_105_501 ();
 FILLCELL_X16 FILLER_105_529 ();
 FILLCELL_X4 FILLER_105_545 ();
 FILLCELL_X1 FILLER_105_576 ();
 FILLCELL_X1 FILLER_105_638 ();
 FILLCELL_X4 FILLER_105_646 ();
 FILLCELL_X2 FILLER_105_650 ();
 FILLCELL_X2 FILLER_105_662 ();
 FILLCELL_X1 FILLER_105_664 ();
 FILLCELL_X1 FILLER_105_668 ();
 FILLCELL_X1 FILLER_105_676 ();
 FILLCELL_X2 FILLER_105_710 ();
 FILLCELL_X4 FILLER_105_721 ();
 FILLCELL_X4 FILLER_105_740 ();
 FILLCELL_X2 FILLER_105_744 ();
 FILLCELL_X4 FILLER_105_779 ();
 FILLCELL_X1 FILLER_105_797 ();
 FILLCELL_X1 FILLER_105_834 ();
 FILLCELL_X1 FILLER_105_844 ();
 FILLCELL_X4 FILLER_105_855 ();
 FILLCELL_X1 FILLER_105_863 ();
 FILLCELL_X1 FILLER_105_870 ();
 FILLCELL_X16 FILLER_105_878 ();
 FILLCELL_X4 FILLER_105_910 ();
 FILLCELL_X2 FILLER_105_914 ();
 FILLCELL_X1 FILLER_105_916 ();
 FILLCELL_X2 FILLER_105_921 ();
 FILLCELL_X4 FILLER_105_927 ();
 FILLCELL_X1 FILLER_105_931 ();
 FILLCELL_X8 FILLER_105_946 ();
 FILLCELL_X4 FILLER_105_954 ();
 FILLCELL_X1 FILLER_105_958 ();
 FILLCELL_X4 FILLER_105_995 ();
 FILLCELL_X1 FILLER_105_999 ();
 FILLCELL_X1 FILLER_105_1037 ();
 FILLCELL_X2 FILLER_105_1058 ();
 FILLCELL_X1 FILLER_105_1060 ();
 FILLCELL_X2 FILLER_105_1078 ();
 FILLCELL_X2 FILLER_105_1089 ();
 FILLCELL_X2 FILLER_105_1115 ();
 FILLCELL_X1 FILLER_105_1117 ();
 FILLCELL_X8 FILLER_105_1125 ();
 FILLCELL_X4 FILLER_105_1133 ();
 FILLCELL_X2 FILLER_105_1144 ();
 FILLCELL_X2 FILLER_105_1155 ();
 FILLCELL_X4 FILLER_105_1179 ();
 FILLCELL_X1 FILLER_105_1183 ();
 FILLCELL_X2 FILLER_105_1187 ();
 FILLCELL_X1 FILLER_105_1189 ();
 FILLCELL_X1 FILLER_105_1207 ();
 FILLCELL_X1 FILLER_105_1245 ();
 FILLCELL_X2 FILLER_105_1252 ();
 FILLCELL_X1 FILLER_105_1254 ();
 FILLCELL_X16 FILLER_106_1 ();
 FILLCELL_X8 FILLER_106_17 ();
 FILLCELL_X4 FILLER_106_25 ();
 FILLCELL_X4 FILLER_106_32 ();
 FILLCELL_X2 FILLER_106_36 ();
 FILLCELL_X1 FILLER_106_38 ();
 FILLCELL_X16 FILLER_106_86 ();
 FILLCELL_X2 FILLER_106_102 ();
 FILLCELL_X1 FILLER_106_156 ();
 FILLCELL_X4 FILLER_106_175 ();
 FILLCELL_X2 FILLER_106_179 ();
 FILLCELL_X1 FILLER_106_181 ();
 FILLCELL_X1 FILLER_106_189 ();
 FILLCELL_X8 FILLER_106_204 ();
 FILLCELL_X2 FILLER_106_212 ();
 FILLCELL_X8 FILLER_106_221 ();
 FILLCELL_X1 FILLER_106_240 ();
 FILLCELL_X2 FILLER_106_245 ();
 FILLCELL_X8 FILLER_106_250 ();
 FILLCELL_X1 FILLER_106_258 ();
 FILLCELL_X2 FILLER_106_263 ();
 FILLCELL_X1 FILLER_106_265 ();
 FILLCELL_X8 FILLER_106_273 ();
 FILLCELL_X4 FILLER_106_281 ();
 FILLCELL_X2 FILLER_106_285 ();
 FILLCELL_X1 FILLER_106_287 ();
 FILLCELL_X4 FILLER_106_308 ();
 FILLCELL_X1 FILLER_106_319 ();
 FILLCELL_X4 FILLER_106_334 ();
 FILLCELL_X2 FILLER_106_338 ();
 FILLCELL_X1 FILLER_106_340 ();
 FILLCELL_X2 FILLER_106_361 ();
 FILLCELL_X1 FILLER_106_363 ();
 FILLCELL_X1 FILLER_106_378 ();
 FILLCELL_X2 FILLER_106_386 ();
 FILLCELL_X1 FILLER_106_388 ();
 FILLCELL_X8 FILLER_106_436 ();
 FILLCELL_X4 FILLER_106_444 ();
 FILLCELL_X4 FILLER_106_462 ();
 FILLCELL_X2 FILLER_106_466 ();
 FILLCELL_X1 FILLER_106_468 ();
 FILLCELL_X2 FILLER_106_476 ();
 FILLCELL_X2 FILLER_106_485 ();
 FILLCELL_X1 FILLER_106_541 ();
 FILLCELL_X1 FILLER_106_549 ();
 FILLCELL_X1 FILLER_106_570 ();
 FILLCELL_X2 FILLER_106_578 ();
 FILLCELL_X2 FILLER_106_587 ();
 FILLCELL_X2 FILLER_106_596 ();
 FILLCELL_X16 FILLER_106_612 ();
 FILLCELL_X2 FILLER_106_628 ();
 FILLCELL_X1 FILLER_106_630 ();
 FILLCELL_X1 FILLER_106_632 ();
 FILLCELL_X8 FILLER_106_640 ();
 FILLCELL_X1 FILLER_106_648 ();
 FILLCELL_X4 FILLER_106_662 ();
 FILLCELL_X1 FILLER_106_666 ();
 FILLCELL_X4 FILLER_106_694 ();
 FILLCELL_X8 FILLER_106_706 ();
 FILLCELL_X4 FILLER_106_714 ();
 FILLCELL_X8 FILLER_106_722 ();
 FILLCELL_X1 FILLER_106_730 ();
 FILLCELL_X1 FILLER_106_776 ();
 FILLCELL_X4 FILLER_106_787 ();
 FILLCELL_X1 FILLER_106_791 ();
 FILLCELL_X8 FILLER_106_799 ();
 FILLCELL_X4 FILLER_106_807 ();
 FILLCELL_X2 FILLER_106_811 ();
 FILLCELL_X2 FILLER_106_856 ();
 FILLCELL_X1 FILLER_106_858 ();
 FILLCELL_X8 FILLER_106_916 ();
 FILLCELL_X1 FILLER_106_924 ();
 FILLCELL_X1 FILLER_106_949 ();
 FILLCELL_X2 FILLER_106_953 ();
 FILLCELL_X1 FILLER_106_955 ();
 FILLCELL_X4 FILLER_106_970 ();
 FILLCELL_X1 FILLER_106_978 ();
 FILLCELL_X8 FILLER_106_989 ();
 FILLCELL_X4 FILLER_106_997 ();
 FILLCELL_X2 FILLER_106_1001 ();
 FILLCELL_X1 FILLER_106_1003 ();
 FILLCELL_X8 FILLER_106_1009 ();
 FILLCELL_X4 FILLER_106_1017 ();
 FILLCELL_X1 FILLER_106_1031 ();
 FILLCELL_X1 FILLER_106_1042 ();
 FILLCELL_X2 FILLER_106_1056 ();
 FILLCELL_X1 FILLER_106_1058 ();
 FILLCELL_X16 FILLER_106_1079 ();
 FILLCELL_X8 FILLER_106_1095 ();
 FILLCELL_X8 FILLER_106_1120 ();
 FILLCELL_X1 FILLER_106_1128 ();
 FILLCELL_X2 FILLER_106_1156 ();
 FILLCELL_X4 FILLER_106_1164 ();
 FILLCELL_X2 FILLER_106_1168 ();
 FILLCELL_X8 FILLER_106_1176 ();
 FILLCELL_X8 FILLER_106_1197 ();
 FILLCELL_X1 FILLER_106_1205 ();
 FILLCELL_X2 FILLER_106_1209 ();
 FILLCELL_X1 FILLER_106_1211 ();
 FILLCELL_X2 FILLER_106_1215 ();
 FILLCELL_X1 FILLER_106_1224 ();
 FILLCELL_X1 FILLER_107_21 ();
 FILLCELL_X1 FILLER_107_50 ();
 FILLCELL_X8 FILLER_107_76 ();
 FILLCELL_X4 FILLER_107_84 ();
 FILLCELL_X2 FILLER_107_88 ();
 FILLCELL_X1 FILLER_107_90 ();
 FILLCELL_X4 FILLER_107_118 ();
 FILLCELL_X2 FILLER_107_122 ();
 FILLCELL_X4 FILLER_107_131 ();
 FILLCELL_X8 FILLER_107_142 ();
 FILLCELL_X1 FILLER_107_150 ();
 FILLCELL_X1 FILLER_107_177 ();
 FILLCELL_X16 FILLER_107_185 ();
 FILLCELL_X2 FILLER_107_221 ();
 FILLCELL_X16 FILLER_107_282 ();
 FILLCELL_X8 FILLER_107_298 ();
 FILLCELL_X1 FILLER_107_306 ();
 FILLCELL_X8 FILLER_107_314 ();
 FILLCELL_X4 FILLER_107_349 ();
 FILLCELL_X2 FILLER_107_353 ();
 FILLCELL_X4 FILLER_107_375 ();
 FILLCELL_X2 FILLER_107_379 ();
 FILLCELL_X1 FILLER_107_401 ();
 FILLCELL_X1 FILLER_107_412 ();
 FILLCELL_X2 FILLER_107_420 ();
 FILLCELL_X1 FILLER_107_422 ();
 FILLCELL_X4 FILLER_107_450 ();
 FILLCELL_X2 FILLER_107_494 ();
 FILLCELL_X16 FILLER_107_501 ();
 FILLCELL_X16 FILLER_107_524 ();
 FILLCELL_X4 FILLER_107_540 ();
 FILLCELL_X2 FILLER_107_544 ();
 FILLCELL_X8 FILLER_107_553 ();
 FILLCELL_X4 FILLER_107_561 ();
 FILLCELL_X2 FILLER_107_565 ();
 FILLCELL_X1 FILLER_107_567 ();
 FILLCELL_X2 FILLER_107_575 ();
 FILLCELL_X2 FILLER_107_584 ();
 FILLCELL_X1 FILLER_107_586 ();
 FILLCELL_X4 FILLER_107_607 ();
 FILLCELL_X1 FILLER_107_611 ();
 FILLCELL_X2 FILLER_107_619 ();
 FILLCELL_X4 FILLER_107_641 ();
 FILLCELL_X1 FILLER_107_645 ();
 FILLCELL_X1 FILLER_107_651 ();
 FILLCELL_X2 FILLER_107_659 ();
 FILLCELL_X8 FILLER_107_686 ();
 FILLCELL_X4 FILLER_107_694 ();
 FILLCELL_X2 FILLER_107_698 ();
 FILLCELL_X1 FILLER_107_700 ();
 FILLCELL_X2 FILLER_107_712 ();
 FILLCELL_X4 FILLER_107_739 ();
 FILLCELL_X2 FILLER_107_743 ();
 FILLCELL_X1 FILLER_107_760 ();
 FILLCELL_X1 FILLER_107_772 ();
 FILLCELL_X4 FILLER_107_784 ();
 FILLCELL_X2 FILLER_107_788 ();
 FILLCELL_X4 FILLER_107_806 ();
 FILLCELL_X1 FILLER_107_810 ();
 FILLCELL_X4 FILLER_107_828 ();
 FILLCELL_X4 FILLER_107_847 ();
 FILLCELL_X1 FILLER_107_851 ();
 FILLCELL_X2 FILLER_107_859 ();
 FILLCELL_X1 FILLER_107_867 ();
 FILLCELL_X1 FILLER_107_874 ();
 FILLCELL_X4 FILLER_107_883 ();
 FILLCELL_X2 FILLER_107_887 ();
 FILLCELL_X1 FILLER_107_889 ();
 FILLCELL_X4 FILLER_107_896 ();
 FILLCELL_X1 FILLER_107_900 ();
 FILLCELL_X4 FILLER_107_912 ();
 FILLCELL_X1 FILLER_107_916 ();
 FILLCELL_X4 FILLER_107_921 ();
 FILLCELL_X2 FILLER_107_925 ();
 FILLCELL_X1 FILLER_107_927 ();
 FILLCELL_X4 FILLER_107_932 ();
 FILLCELL_X2 FILLER_107_936 ();
 FILLCELL_X1 FILLER_107_938 ();
 FILLCELL_X1 FILLER_107_959 ();
 FILLCELL_X16 FILLER_107_979 ();
 FILLCELL_X8 FILLER_107_995 ();
 FILLCELL_X1 FILLER_107_1003 ();
 FILLCELL_X1 FILLER_107_1009 ();
 FILLCELL_X1 FILLER_107_1025 ();
 FILLCELL_X2 FILLER_107_1036 ();
 FILLCELL_X1 FILLER_107_1038 ();
 FILLCELL_X2 FILLER_107_1067 ();
 FILLCELL_X1 FILLER_107_1075 ();
 FILLCELL_X1 FILLER_107_1086 ();
 FILLCELL_X1 FILLER_107_1089 ();
 FILLCELL_X16 FILLER_107_1099 ();
 FILLCELL_X8 FILLER_107_1115 ();
 FILLCELL_X1 FILLER_107_1123 ();
 FILLCELL_X8 FILLER_107_1137 ();
 FILLCELL_X2 FILLER_107_1145 ();
 FILLCELL_X2 FILLER_107_1154 ();
 FILLCELL_X1 FILLER_107_1156 ();
 FILLCELL_X2 FILLER_107_1189 ();
 FILLCELL_X4 FILLER_107_1196 ();
 FILLCELL_X1 FILLER_107_1200 ();
 FILLCELL_X2 FILLER_107_1207 ();
 FILLCELL_X1 FILLER_107_1209 ();
 FILLCELL_X2 FILLER_107_1250 ();
 FILLCELL_X8 FILLER_108_1 ();
 FILLCELL_X4 FILLER_108_9 ();
 FILLCELL_X4 FILLER_108_27 ();
 FILLCELL_X2 FILLER_108_31 ();
 FILLCELL_X2 FILLER_108_40 ();
 FILLCELL_X4 FILLER_108_62 ();
 FILLCELL_X2 FILLER_108_66 ();
 FILLCELL_X4 FILLER_108_89 ();
 FILLCELL_X2 FILLER_108_93 ();
 FILLCELL_X8 FILLER_108_102 ();
 FILLCELL_X2 FILLER_108_110 ();
 FILLCELL_X1 FILLER_108_126 ();
 FILLCELL_X1 FILLER_108_174 ();
 FILLCELL_X1 FILLER_108_179 ();
 FILLCELL_X1 FILLER_108_186 ();
 FILLCELL_X1 FILLER_108_201 ();
 FILLCELL_X1 FILLER_108_222 ();
 FILLCELL_X1 FILLER_108_243 ();
 FILLCELL_X1 FILLER_108_248 ();
 FILLCELL_X2 FILLER_108_252 ();
 FILLCELL_X2 FILLER_108_271 ();
 FILLCELL_X4 FILLER_108_294 ();
 FILLCELL_X2 FILLER_108_298 ();
 FILLCELL_X1 FILLER_108_300 ();
 FILLCELL_X4 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_332 ();
 FILLCELL_X2 FILLER_108_364 ();
 FILLCELL_X1 FILLER_108_366 ();
 FILLCELL_X16 FILLER_108_374 ();
 FILLCELL_X1 FILLER_108_390 ();
 FILLCELL_X1 FILLER_108_409 ();
 FILLCELL_X2 FILLER_108_433 ();
 FILLCELL_X2 FILLER_108_442 ();
 FILLCELL_X1 FILLER_108_444 ();
 FILLCELL_X2 FILLER_108_452 ();
 FILLCELL_X2 FILLER_108_461 ();
 FILLCELL_X2 FILLER_108_470 ();
 FILLCELL_X1 FILLER_108_472 ();
 FILLCELL_X4 FILLER_108_480 ();
 FILLCELL_X1 FILLER_108_484 ();
 FILLCELL_X4 FILLER_108_492 ();
 FILLCELL_X1 FILLER_108_496 ();
 FILLCELL_X4 FILLER_108_500 ();
 FILLCELL_X1 FILLER_108_518 ();
 FILLCELL_X2 FILLER_108_526 ();
 FILLCELL_X1 FILLER_108_548 ();
 FILLCELL_X2 FILLER_108_569 ();
 FILLCELL_X16 FILLER_108_591 ();
 FILLCELL_X4 FILLER_108_607 ();
 FILLCELL_X1 FILLER_108_611 ();
 FILLCELL_X8 FILLER_108_619 ();
 FILLCELL_X4 FILLER_108_627 ();
 FILLCELL_X16 FILLER_108_642 ();
 FILLCELL_X8 FILLER_108_658 ();
 FILLCELL_X4 FILLER_108_666 ();
 FILLCELL_X1 FILLER_108_670 ();
 FILLCELL_X1 FILLER_108_675 ();
 FILLCELL_X1 FILLER_108_700 ();
 FILLCELL_X4 FILLER_108_712 ();
 FILLCELL_X2 FILLER_108_716 ();
 FILLCELL_X2 FILLER_108_729 ();
 FILLCELL_X1 FILLER_108_736 ();
 FILLCELL_X2 FILLER_108_753 ();
 FILLCELL_X1 FILLER_108_755 ();
 FILLCELL_X2 FILLER_108_758 ();
 FILLCELL_X8 FILLER_108_769 ();
 FILLCELL_X1 FILLER_108_796 ();
 FILLCELL_X1 FILLER_108_804 ();
 FILLCELL_X4 FILLER_108_812 ();
 FILLCELL_X2 FILLER_108_822 ();
 FILLCELL_X1 FILLER_108_824 ();
 FILLCELL_X1 FILLER_108_831 ();
 FILLCELL_X1 FILLER_108_846 ();
 FILLCELL_X2 FILLER_108_854 ();
 FILLCELL_X1 FILLER_108_856 ();
 FILLCELL_X1 FILLER_108_863 ();
 FILLCELL_X4 FILLER_108_871 ();
 FILLCELL_X1 FILLER_108_875 ();
 FILLCELL_X2 FILLER_108_886 ();
 FILLCELL_X1 FILLER_108_888 ();
 FILLCELL_X2 FILLER_108_899 ();
 FILLCELL_X4 FILLER_108_915 ();
 FILLCELL_X2 FILLER_108_919 ();
 FILLCELL_X1 FILLER_108_921 ();
 FILLCELL_X1 FILLER_108_926 ();
 FILLCELL_X2 FILLER_108_944 ();
 FILLCELL_X1 FILLER_108_946 ();
 FILLCELL_X2 FILLER_108_967 ();
 FILLCELL_X4 FILLER_108_986 ();
 FILLCELL_X2 FILLER_108_990 ();
 FILLCELL_X1 FILLER_108_992 ();
 FILLCELL_X4 FILLER_108_997 ();
 FILLCELL_X1 FILLER_108_1001 ();
 FILLCELL_X4 FILLER_108_1017 ();
 FILLCELL_X1 FILLER_108_1021 ();
 FILLCELL_X1 FILLER_108_1029 ();
 FILLCELL_X2 FILLER_108_1035 ();
 FILLCELL_X1 FILLER_108_1051 ();
 FILLCELL_X1 FILLER_108_1062 ();
 FILLCELL_X1 FILLER_108_1079 ();
 FILLCELL_X1 FILLER_108_1088 ();
 FILLCELL_X1 FILLER_108_1096 ();
 FILLCELL_X1 FILLER_108_1101 ();
 FILLCELL_X2 FILLER_108_1109 ();
 FILLCELL_X4 FILLER_108_1135 ();
 FILLCELL_X1 FILLER_108_1139 ();
 FILLCELL_X2 FILLER_108_1148 ();
 FILLCELL_X4 FILLER_108_1168 ();
 FILLCELL_X1 FILLER_108_1172 ();
 FILLCELL_X1 FILLER_108_1179 ();
 FILLCELL_X8 FILLER_108_1214 ();
 FILLCELL_X1 FILLER_108_1222 ();
 FILLCELL_X4 FILLER_108_1228 ();
 FILLCELL_X2 FILLER_108_1232 ();
 FILLCELL_X2 FILLER_108_1250 ();
 FILLCELL_X2 FILLER_109_1 ();
 FILLCELL_X4 FILLER_109_23 ();
 FILLCELL_X2 FILLER_109_27 ();
 FILLCELL_X4 FILLER_109_50 ();
 FILLCELL_X16 FILLER_109_82 ();
 FILLCELL_X4 FILLER_109_98 ();
 FILLCELL_X2 FILLER_109_102 ();
 FILLCELL_X32 FILLER_109_139 ();
 FILLCELL_X4 FILLER_109_171 ();
 FILLCELL_X2 FILLER_109_175 ();
 FILLCELL_X4 FILLER_109_182 ();
 FILLCELL_X2 FILLER_109_238 ();
 FILLCELL_X4 FILLER_109_260 ();
 FILLCELL_X2 FILLER_109_264 ();
 FILLCELL_X4 FILLER_109_273 ();
 FILLCELL_X2 FILLER_109_277 ();
 FILLCELL_X4 FILLER_109_296 ();
 FILLCELL_X2 FILLER_109_300 ();
 FILLCELL_X1 FILLER_109_302 ();
 FILLCELL_X4 FILLER_109_307 ();
 FILLCELL_X2 FILLER_109_320 ();
 FILLCELL_X2 FILLER_109_328 ();
 FILLCELL_X1 FILLER_109_407 ();
 FILLCELL_X4 FILLER_109_422 ();
 FILLCELL_X1 FILLER_109_426 ();
 FILLCELL_X8 FILLER_109_470 ();
 FILLCELL_X4 FILLER_109_478 ();
 FILLCELL_X1 FILLER_109_482 ();
 FILLCELL_X8 FILLER_109_504 ();
 FILLCELL_X4 FILLER_109_512 ();
 FILLCELL_X2 FILLER_109_530 ();
 FILLCELL_X16 FILLER_109_539 ();
 FILLCELL_X2 FILLER_109_555 ();
 FILLCELL_X4 FILLER_109_561 ();
 FILLCELL_X2 FILLER_109_565 ();
 FILLCELL_X1 FILLER_109_567 ();
 FILLCELL_X4 FILLER_109_575 ();
 FILLCELL_X1 FILLER_109_579 ();
 FILLCELL_X1 FILLER_109_593 ();
 FILLCELL_X1 FILLER_109_602 ();
 FILLCELL_X4 FILLER_109_610 ();
 FILLCELL_X2 FILLER_109_614 ();
 FILLCELL_X8 FILLER_109_636 ();
 FILLCELL_X4 FILLER_109_644 ();
 FILLCELL_X2 FILLER_109_648 ();
 FILLCELL_X16 FILLER_109_655 ();
 FILLCELL_X8 FILLER_109_671 ();
 FILLCELL_X2 FILLER_109_679 ();
 FILLCELL_X2 FILLER_109_686 ();
 FILLCELL_X1 FILLER_109_688 ();
 FILLCELL_X4 FILLER_109_702 ();
 FILLCELL_X2 FILLER_109_706 ();
 FILLCELL_X4 FILLER_109_723 ();
 FILLCELL_X1 FILLER_109_760 ();
 FILLCELL_X4 FILLER_109_771 ();
 FILLCELL_X1 FILLER_109_775 ();
 FILLCELL_X1 FILLER_109_790 ();
 FILLCELL_X2 FILLER_109_803 ();
 FILLCELL_X4 FILLER_109_825 ();
 FILLCELL_X2 FILLER_109_829 ();
 FILLCELL_X1 FILLER_109_831 ();
 FILLCELL_X1 FILLER_109_839 ();
 FILLCELL_X1 FILLER_109_852 ();
 FILLCELL_X1 FILLER_109_860 ();
 FILLCELL_X1 FILLER_109_871 ();
 FILLCELL_X2 FILLER_109_882 ();
 FILLCELL_X1 FILLER_109_884 ();
 FILLCELL_X1 FILLER_109_904 ();
 FILLCELL_X2 FILLER_109_909 ();
 FILLCELL_X1 FILLER_109_911 ();
 FILLCELL_X8 FILLER_109_940 ();
 FILLCELL_X4 FILLER_109_948 ();
 FILLCELL_X1 FILLER_109_952 ();
 FILLCELL_X1 FILLER_109_963 ();
 FILLCELL_X8 FILLER_109_984 ();
 FILLCELL_X4 FILLER_109_992 ();
 FILLCELL_X1 FILLER_109_996 ();
 FILLCELL_X4 FILLER_109_1009 ();
 FILLCELL_X1 FILLER_109_1028 ();
 FILLCELL_X8 FILLER_109_1033 ();
 FILLCELL_X1 FILLER_109_1041 ();
 FILLCELL_X1 FILLER_109_1051 ();
 FILLCELL_X4 FILLER_109_1055 ();
 FILLCELL_X1 FILLER_109_1059 ();
 FILLCELL_X2 FILLER_109_1071 ();
 FILLCELL_X1 FILLER_109_1077 ();
 FILLCELL_X8 FILLER_109_1090 ();
 FILLCELL_X1 FILLER_109_1098 ();
 FILLCELL_X2 FILLER_109_1107 ();
 FILLCELL_X8 FILLER_109_1116 ();
 FILLCELL_X4 FILLER_109_1124 ();
 FILLCELL_X2 FILLER_109_1128 ();
 FILLCELL_X32 FILLER_109_1136 ();
 FILLCELL_X4 FILLER_109_1168 ();
 FILLCELL_X1 FILLER_109_1174 ();
 FILLCELL_X4 FILLER_109_1185 ();
 FILLCELL_X1 FILLER_109_1189 ();
 FILLCELL_X4 FILLER_109_1201 ();
 FILLCELL_X2 FILLER_109_1224 ();
 FILLCELL_X8 FILLER_110_1 ();
 FILLCELL_X4 FILLER_110_9 ();
 FILLCELL_X1 FILLER_110_13 ();
 FILLCELL_X2 FILLER_110_41 ();
 FILLCELL_X1 FILLER_110_66 ();
 FILLCELL_X1 FILLER_110_108 ();
 FILLCELL_X1 FILLER_110_116 ();
 FILLCELL_X1 FILLER_110_124 ();
 FILLCELL_X2 FILLER_110_166 ();
 FILLCELL_X1 FILLER_110_179 ();
 FILLCELL_X8 FILLER_110_184 ();
 FILLCELL_X1 FILLER_110_192 ();
 FILLCELL_X1 FILLER_110_216 ();
 FILLCELL_X2 FILLER_110_224 ();
 FILLCELL_X2 FILLER_110_233 ();
 FILLCELL_X8 FILLER_110_255 ();
 FILLCELL_X1 FILLER_110_263 ();
 FILLCELL_X2 FILLER_110_302 ();
 FILLCELL_X1 FILLER_110_307 ();
 FILLCELL_X2 FILLER_110_328 ();
 FILLCELL_X1 FILLER_110_330 ();
 FILLCELL_X4 FILLER_110_358 ();
 FILLCELL_X2 FILLER_110_362 ();
 FILLCELL_X1 FILLER_110_364 ();
 FILLCELL_X4 FILLER_110_379 ();
 FILLCELL_X2 FILLER_110_383 ();
 FILLCELL_X4 FILLER_110_392 ();
 FILLCELL_X4 FILLER_110_399 ();
 FILLCELL_X2 FILLER_110_403 ();
 FILLCELL_X1 FILLER_110_405 ();
 FILLCELL_X1 FILLER_110_410 ();
 FILLCELL_X2 FILLER_110_414 ();
 FILLCELL_X1 FILLER_110_416 ();
 FILLCELL_X4 FILLER_110_424 ();
 FILLCELL_X16 FILLER_110_438 ();
 FILLCELL_X8 FILLER_110_454 ();
 FILLCELL_X1 FILLER_110_465 ();
 FILLCELL_X2 FILLER_110_486 ();
 FILLCELL_X1 FILLER_110_488 ();
 FILLCELL_X2 FILLER_110_496 ();
 FILLCELL_X2 FILLER_110_510 ();
 FILLCELL_X1 FILLER_110_512 ();
 FILLCELL_X4 FILLER_110_525 ();
 FILLCELL_X4 FILLER_110_536 ();
 FILLCELL_X1 FILLER_110_540 ();
 FILLCELL_X8 FILLER_110_548 ();
 FILLCELL_X2 FILLER_110_556 ();
 FILLCELL_X1 FILLER_110_558 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_639 ();
 FILLCELL_X16 FILLER_110_671 ();
 FILLCELL_X4 FILLER_110_687 ();
 FILLCELL_X2 FILLER_110_746 ();
 FILLCELL_X1 FILLER_110_748 ();
 FILLCELL_X8 FILLER_110_772 ();
 FILLCELL_X4 FILLER_110_780 ();
 FILLCELL_X16 FILLER_110_791 ();
 FILLCELL_X8 FILLER_110_807 ();
 FILLCELL_X4 FILLER_110_822 ();
 FILLCELL_X2 FILLER_110_826 ();
 FILLCELL_X4 FILLER_110_831 ();
 FILLCELL_X2 FILLER_110_846 ();
 FILLCELL_X1 FILLER_110_848 ();
 FILLCELL_X4 FILLER_110_855 ();
 FILLCELL_X1 FILLER_110_859 ();
 FILLCELL_X8 FILLER_110_874 ();
 FILLCELL_X4 FILLER_110_882 ();
 FILLCELL_X2 FILLER_110_891 ();
 FILLCELL_X1 FILLER_110_893 ();
 FILLCELL_X4 FILLER_110_901 ();
 FILLCELL_X2 FILLER_110_905 ();
 FILLCELL_X8 FILLER_110_914 ();
 FILLCELL_X2 FILLER_110_922 ();
 FILLCELL_X1 FILLER_110_924 ();
 FILLCELL_X4 FILLER_110_929 ();
 FILLCELL_X2 FILLER_110_933 ();
 FILLCELL_X1 FILLER_110_935 ();
 FILLCELL_X1 FILLER_110_950 ();
 FILLCELL_X2 FILLER_110_959 ();
 FILLCELL_X2 FILLER_110_979 ();
 FILLCELL_X8 FILLER_110_995 ();
 FILLCELL_X2 FILLER_110_1003 ();
 FILLCELL_X1 FILLER_110_1028 ();
 FILLCELL_X4 FILLER_110_1036 ();
 FILLCELL_X1 FILLER_110_1040 ();
 FILLCELL_X2 FILLER_110_1045 ();
 FILLCELL_X2 FILLER_110_1058 ();
 FILLCELL_X1 FILLER_110_1060 ();
 FILLCELL_X4 FILLER_110_1072 ();
 FILLCELL_X1 FILLER_110_1076 ();
 FILLCELL_X2 FILLER_110_1087 ();
 FILLCELL_X4 FILLER_110_1091 ();
 FILLCELL_X1 FILLER_110_1095 ();
 FILLCELL_X4 FILLER_110_1121 ();
 FILLCELL_X2 FILLER_110_1125 ();
 FILLCELL_X1 FILLER_110_1127 ();
 FILLCELL_X2 FILLER_110_1152 ();
 FILLCELL_X8 FILLER_110_1200 ();
 FILLCELL_X2 FILLER_110_1208 ();
 FILLCELL_X1 FILLER_110_1225 ();
 FILLCELL_X8 FILLER_110_1231 ();
 FILLCELL_X4 FILLER_110_1239 ();
 FILLCELL_X2 FILLER_110_1249 ();
 FILLCELL_X1 FILLER_110_1251 ();
 FILLCELL_X2 FILLER_111_28 ();
 FILLCELL_X4 FILLER_111_37 ();
 FILLCELL_X1 FILLER_111_41 ();
 FILLCELL_X4 FILLER_111_83 ();
 FILLCELL_X4 FILLER_111_114 ();
 FILLCELL_X2 FILLER_111_118 ();
 FILLCELL_X16 FILLER_111_140 ();
 FILLCELL_X2 FILLER_111_156 ();
 FILLCELL_X2 FILLER_111_179 ();
 FILLCELL_X2 FILLER_111_192 ();
 FILLCELL_X1 FILLER_111_194 ();
 FILLCELL_X1 FILLER_111_209 ();
 FILLCELL_X2 FILLER_111_242 ();
 FILLCELL_X16 FILLER_111_247 ();
 FILLCELL_X2 FILLER_111_263 ();
 FILLCELL_X4 FILLER_111_268 ();
 FILLCELL_X2 FILLER_111_272 ();
 FILLCELL_X8 FILLER_111_281 ();
 FILLCELL_X4 FILLER_111_289 ();
 FILLCELL_X2 FILLER_111_313 ();
 FILLCELL_X4 FILLER_111_329 ();
 FILLCELL_X1 FILLER_111_333 ();
 FILLCELL_X16 FILLER_111_337 ();
 FILLCELL_X8 FILLER_111_353 ();
 FILLCELL_X1 FILLER_111_361 ();
 FILLCELL_X8 FILLER_111_376 ();
 FILLCELL_X4 FILLER_111_411 ();
 FILLCELL_X2 FILLER_111_415 ();
 FILLCELL_X4 FILLER_111_421 ();
 FILLCELL_X1 FILLER_111_425 ();
 FILLCELL_X2 FILLER_111_446 ();
 FILLCELL_X4 FILLER_111_461 ();
 FILLCELL_X2 FILLER_111_465 ();
 FILLCELL_X4 FILLER_111_499 ();
 FILLCELL_X2 FILLER_111_503 ();
 FILLCELL_X1 FILLER_111_512 ();
 FILLCELL_X8 FILLER_111_601 ();
 FILLCELL_X4 FILLER_111_609 ();
 FILLCELL_X4 FILLER_111_627 ();
 FILLCELL_X1 FILLER_111_631 ();
 FILLCELL_X2 FILLER_111_649 ();
 FILLCELL_X1 FILLER_111_651 ();
 FILLCELL_X1 FILLER_111_659 ();
 FILLCELL_X16 FILLER_111_687 ();
 FILLCELL_X8 FILLER_111_703 ();
 FILLCELL_X2 FILLER_111_711 ();
 FILLCELL_X1 FILLER_111_723 ();
 FILLCELL_X2 FILLER_111_733 ();
 FILLCELL_X2 FILLER_111_740 ();
 FILLCELL_X2 FILLER_111_755 ();
 FILLCELL_X1 FILLER_111_757 ();
 FILLCELL_X8 FILLER_111_767 ();
 FILLCELL_X1 FILLER_111_775 ();
 FILLCELL_X4 FILLER_111_793 ();
 FILLCELL_X2 FILLER_111_804 ();
 FILLCELL_X1 FILLER_111_806 ();
 FILLCELL_X4 FILLER_111_814 ();
 FILLCELL_X1 FILLER_111_831 ();
 FILLCELL_X1 FILLER_111_845 ();
 FILLCELL_X1 FILLER_111_850 ();
 FILLCELL_X4 FILLER_111_858 ();
 FILLCELL_X2 FILLER_111_862 ();
 FILLCELL_X1 FILLER_111_864 ();
 FILLCELL_X4 FILLER_111_872 ();
 FILLCELL_X2 FILLER_111_876 ();
 FILLCELL_X8 FILLER_111_893 ();
 FILLCELL_X2 FILLER_111_901 ();
 FILLCELL_X1 FILLER_111_903 ();
 FILLCELL_X4 FILLER_111_909 ();
 FILLCELL_X2 FILLER_111_913 ();
 FILLCELL_X1 FILLER_111_915 ();
 FILLCELL_X2 FILLER_111_931 ();
 FILLCELL_X1 FILLER_111_933 ();
 FILLCELL_X1 FILLER_111_936 ();
 FILLCELL_X8 FILLER_111_942 ();
 FILLCELL_X4 FILLER_111_955 ();
 FILLCELL_X2 FILLER_111_1027 ();
 FILLCELL_X4 FILLER_111_1043 ();
 FILLCELL_X2 FILLER_111_1047 ();
 FILLCELL_X1 FILLER_111_1064 ();
 FILLCELL_X1 FILLER_111_1069 ();
 FILLCELL_X2 FILLER_111_1074 ();
 FILLCELL_X2 FILLER_111_1083 ();
 FILLCELL_X2 FILLER_111_1104 ();
 FILLCELL_X8 FILLER_111_1109 ();
 FILLCELL_X1 FILLER_111_1117 ();
 FILLCELL_X4 FILLER_111_1135 ();
 FILLCELL_X8 FILLER_111_1156 ();
 FILLCELL_X1 FILLER_111_1164 ();
 FILLCELL_X8 FILLER_111_1201 ();
 FILLCELL_X4 FILLER_111_1209 ();
 FILLCELL_X4 FILLER_111_1217 ();
 FILLCELL_X4 FILLER_111_1228 ();
 FILLCELL_X1 FILLER_111_1232 ();
 FILLCELL_X4 FILLER_111_1236 ();
 FILLCELL_X2 FILLER_111_1240 ();
 FILLCELL_X1 FILLER_111_1242 ();
 FILLCELL_X1 FILLER_111_1246 ();
 FILLCELL_X2 FILLER_111_1253 ();
 FILLCELL_X8 FILLER_112_1 ();
 FILLCELL_X4 FILLER_112_9 ();
 FILLCELL_X1 FILLER_112_13 ();
 FILLCELL_X8 FILLER_112_19 ();
 FILLCELL_X2 FILLER_112_27 ();
 FILLCELL_X16 FILLER_112_43 ();
 FILLCELL_X8 FILLER_112_59 ();
 FILLCELL_X1 FILLER_112_81 ();
 FILLCELL_X16 FILLER_112_89 ();
 FILLCELL_X8 FILLER_112_105 ();
 FILLCELL_X2 FILLER_112_125 ();
 FILLCELL_X4 FILLER_112_168 ();
 FILLCELL_X2 FILLER_112_172 ();
 FILLCELL_X8 FILLER_112_181 ();
 FILLCELL_X4 FILLER_112_189 ();
 FILLCELL_X2 FILLER_112_193 ();
 FILLCELL_X1 FILLER_112_195 ();
 FILLCELL_X1 FILLER_112_231 ();
 FILLCELL_X1 FILLER_112_279 ();
 FILLCELL_X4 FILLER_112_287 ();
 FILLCELL_X2 FILLER_112_298 ();
 FILLCELL_X4 FILLER_112_307 ();
 FILLCELL_X2 FILLER_112_311 ();
 FILLCELL_X1 FILLER_112_334 ();
 FILLCELL_X8 FILLER_112_362 ();
 FILLCELL_X2 FILLER_112_370 ();
 FILLCELL_X32 FILLER_112_379 ();
 FILLCELL_X1 FILLER_112_411 ();
 FILLCELL_X8 FILLER_112_419 ();
 FILLCELL_X2 FILLER_112_427 ();
 FILLCELL_X1 FILLER_112_449 ();
 FILLCELL_X2 FILLER_112_492 ();
 FILLCELL_X2 FILLER_112_521 ();
 FILLCELL_X16 FILLER_112_543 ();
 FILLCELL_X4 FILLER_112_570 ();
 FILLCELL_X2 FILLER_112_574 ();
 FILLCELL_X1 FILLER_112_576 ();
 FILLCELL_X8 FILLER_112_632 ();
 FILLCELL_X4 FILLER_112_640 ();
 FILLCELL_X2 FILLER_112_644 ();
 FILLCELL_X4 FILLER_112_650 ();
 FILLCELL_X2 FILLER_112_654 ();
 FILLCELL_X1 FILLER_112_656 ();
 FILLCELL_X1 FILLER_112_671 ();
 FILLCELL_X2 FILLER_112_682 ();
 FILLCELL_X1 FILLER_112_684 ();
 FILLCELL_X2 FILLER_112_712 ();
 FILLCELL_X4 FILLER_112_734 ();
 FILLCELL_X4 FILLER_112_748 ();
 FILLCELL_X2 FILLER_112_752 ();
 FILLCELL_X1 FILLER_112_754 ();
 FILLCELL_X8 FILLER_112_762 ();
 FILLCELL_X2 FILLER_112_770 ();
 FILLCELL_X1 FILLER_112_780 ();
 FILLCELL_X1 FILLER_112_785 ();
 FILLCELL_X1 FILLER_112_790 ();
 FILLCELL_X1 FILLER_112_807 ();
 FILLCELL_X1 FILLER_112_812 ();
 FILLCELL_X8 FILLER_112_821 ();
 FILLCELL_X1 FILLER_112_829 ();
 FILLCELL_X16 FILLER_112_844 ();
 FILLCELL_X2 FILLER_112_860 ();
 FILLCELL_X2 FILLER_112_877 ();
 FILLCELL_X4 FILLER_112_889 ();
 FILLCELL_X4 FILLER_112_913 ();
 FILLCELL_X2 FILLER_112_922 ();
 FILLCELL_X4 FILLER_112_929 ();
 FILLCELL_X2 FILLER_112_933 ();
 FILLCELL_X8 FILLER_112_959 ();
 FILLCELL_X4 FILLER_112_967 ();
 FILLCELL_X2 FILLER_112_971 ();
 FILLCELL_X16 FILLER_112_988 ();
 FILLCELL_X8 FILLER_112_1004 ();
 FILLCELL_X1 FILLER_112_1012 ();
 FILLCELL_X2 FILLER_112_1053 ();
 FILLCELL_X1 FILLER_112_1055 ();
 FILLCELL_X16 FILLER_112_1087 ();
 FILLCELL_X8 FILLER_112_1103 ();
 FILLCELL_X4 FILLER_112_1111 ();
 FILLCELL_X2 FILLER_112_1115 ();
 FILLCELL_X1 FILLER_112_1117 ();
 FILLCELL_X4 FILLER_112_1137 ();
 FILLCELL_X2 FILLER_112_1141 ();
 FILLCELL_X1 FILLER_112_1150 ();
 FILLCELL_X2 FILLER_112_1198 ();
 FILLCELL_X1 FILLER_112_1220 ();
 FILLCELL_X16 FILLER_112_1231 ();
 FILLCELL_X8 FILLER_112_1247 ();
 FILLCELL_X2 FILLER_113_1 ();
 FILLCELL_X8 FILLER_113_37 ();
 FILLCELL_X4 FILLER_113_45 ();
 FILLCELL_X2 FILLER_113_49 ();
 FILLCELL_X1 FILLER_113_51 ();
 FILLCELL_X4 FILLER_113_59 ();
 FILLCELL_X2 FILLER_113_63 ();
 FILLCELL_X2 FILLER_113_85 ();
 FILLCELL_X8 FILLER_113_114 ();
 FILLCELL_X2 FILLER_113_122 ();
 FILLCELL_X1 FILLER_113_124 ();
 FILLCELL_X2 FILLER_113_172 ();
 FILLCELL_X1 FILLER_113_174 ();
 FILLCELL_X4 FILLER_113_216 ();
 FILLCELL_X2 FILLER_113_220 ();
 FILLCELL_X1 FILLER_113_222 ();
 FILLCELL_X4 FILLER_113_227 ();
 FILLCELL_X2 FILLER_113_231 ();
 FILLCELL_X1 FILLER_113_233 ();
 FILLCELL_X1 FILLER_113_237 ();
 FILLCELL_X4 FILLER_113_245 ();
 FILLCELL_X1 FILLER_113_253 ();
 FILLCELL_X4 FILLER_113_257 ();
 FILLCELL_X8 FILLER_113_286 ();
 FILLCELL_X1 FILLER_113_294 ();
 FILLCELL_X4 FILLER_113_315 ();
 FILLCELL_X4 FILLER_113_326 ();
 FILLCELL_X2 FILLER_113_330 ();
 FILLCELL_X1 FILLER_113_332 ();
 FILLCELL_X4 FILLER_113_353 ();
 FILLCELL_X1 FILLER_113_357 ();
 FILLCELL_X4 FILLER_113_414 ();
 FILLCELL_X2 FILLER_113_418 ();
 FILLCELL_X4 FILLER_113_438 ();
 FILLCELL_X1 FILLER_113_442 ();
 FILLCELL_X4 FILLER_113_500 ();
 FILLCELL_X4 FILLER_113_545 ();
 FILLCELL_X1 FILLER_113_557 ();
 FILLCELL_X2 FILLER_113_590 ();
 FILLCELL_X8 FILLER_113_599 ();
 FILLCELL_X1 FILLER_113_607 ();
 FILLCELL_X2 FILLER_113_615 ();
 FILLCELL_X1 FILLER_113_617 ();
 FILLCELL_X1 FILLER_113_632 ();
 FILLCELL_X8 FILLER_113_650 ();
 FILLCELL_X4 FILLER_113_658 ();
 FILLCELL_X1 FILLER_113_662 ();
 FILLCELL_X2 FILLER_113_695 ();
 FILLCELL_X1 FILLER_113_697 ();
 FILLCELL_X2 FILLER_113_704 ();
 FILLCELL_X1 FILLER_113_709 ();
 FILLCELL_X4 FILLER_113_737 ();
 FILLCELL_X4 FILLER_113_749 ();
 FILLCELL_X4 FILLER_113_757 ();
 FILLCELL_X4 FILLER_113_765 ();
 FILLCELL_X8 FILLER_113_772 ();
 FILLCELL_X1 FILLER_113_787 ();
 FILLCELL_X2 FILLER_113_795 ();
 FILLCELL_X1 FILLER_113_797 ();
 FILLCELL_X1 FILLER_113_817 ();
 FILLCELL_X8 FILLER_113_821 ();
 FILLCELL_X4 FILLER_113_829 ();
 FILLCELL_X16 FILLER_113_840 ();
 FILLCELL_X1 FILLER_113_856 ();
 FILLCELL_X8 FILLER_113_865 ();
 FILLCELL_X4 FILLER_113_873 ();
 FILLCELL_X1 FILLER_113_877 ();
 FILLCELL_X4 FILLER_113_882 ();
 FILLCELL_X2 FILLER_113_886 ();
 FILLCELL_X1 FILLER_113_895 ();
 FILLCELL_X1 FILLER_113_905 ();
 FILLCELL_X4 FILLER_113_911 ();
 FILLCELL_X2 FILLER_113_915 ();
 FILLCELL_X2 FILLER_113_927 ();
 FILLCELL_X2 FILLER_113_934 ();
 FILLCELL_X1 FILLER_113_936 ();
 FILLCELL_X8 FILLER_113_947 ();
 FILLCELL_X4 FILLER_113_955 ();
 FILLCELL_X1 FILLER_113_981 ();
 FILLCELL_X4 FILLER_113_1004 ();
 FILLCELL_X1 FILLER_113_1030 ();
 FILLCELL_X8 FILLER_113_1047 ();
 FILLCELL_X4 FILLER_113_1055 ();
 FILLCELL_X2 FILLER_113_1059 ();
 FILLCELL_X8 FILLER_113_1086 ();
 FILLCELL_X4 FILLER_113_1094 ();
 FILLCELL_X1 FILLER_113_1098 ();
 FILLCELL_X2 FILLER_113_1133 ();
 FILLCELL_X4 FILLER_113_1159 ();
 FILLCELL_X2 FILLER_113_1163 ();
 FILLCELL_X1 FILLER_113_1165 ();
 FILLCELL_X4 FILLER_113_1202 ();
 FILLCELL_X1 FILLER_113_1216 ();
 FILLCELL_X2 FILLER_113_1234 ();
 FILLCELL_X1 FILLER_113_1236 ();
 FILLCELL_X4 FILLER_113_1240 ();
 FILLCELL_X2 FILLER_113_1244 ();
 FILLCELL_X4 FILLER_113_1249 ();
 FILLCELL_X2 FILLER_113_1253 ();
 FILLCELL_X4 FILLER_114_21 ();
 FILLCELL_X1 FILLER_114_39 ();
 FILLCELL_X1 FILLER_114_87 ();
 FILLCELL_X2 FILLER_114_133 ();
 FILLCELL_X1 FILLER_114_135 ();
 FILLCELL_X4 FILLER_114_143 ();
 FILLCELL_X2 FILLER_114_147 ();
 FILLCELL_X1 FILLER_114_149 ();
 FILLCELL_X2 FILLER_114_162 ();
 FILLCELL_X1 FILLER_114_164 ();
 FILLCELL_X2 FILLER_114_179 ();
 FILLCELL_X8 FILLER_114_188 ();
 FILLCELL_X1 FILLER_114_196 ();
 FILLCELL_X2 FILLER_114_237 ();
 FILLCELL_X4 FILLER_114_279 ();
 FILLCELL_X8 FILLER_114_287 ();
 FILLCELL_X8 FILLER_114_298 ();
 FILLCELL_X2 FILLER_114_306 ();
 FILLCELL_X1 FILLER_114_308 ();
 FILLCELL_X4 FILLER_114_329 ();
 FILLCELL_X1 FILLER_114_333 ();
 FILLCELL_X2 FILLER_114_341 ();
 FILLCELL_X1 FILLER_114_343 ();
 FILLCELL_X8 FILLER_114_364 ();
 FILLCELL_X4 FILLER_114_372 ();
 FILLCELL_X1 FILLER_114_376 ();
 FILLCELL_X4 FILLER_114_398 ();
 FILLCELL_X1 FILLER_114_438 ();
 FILLCELL_X1 FILLER_114_442 ();
 FILLCELL_X1 FILLER_114_450 ();
 FILLCELL_X1 FILLER_114_458 ();
 FILLCELL_X4 FILLER_114_522 ();
 FILLCELL_X1 FILLER_114_526 ();
 FILLCELL_X4 FILLER_114_531 ();
 FILLCELL_X1 FILLER_114_535 ();
 FILLCELL_X32 FILLER_114_543 ();
 FILLCELL_X2 FILLER_114_575 ();
 FILLCELL_X1 FILLER_114_577 ();
 FILLCELL_X8 FILLER_114_592 ();
 FILLCELL_X2 FILLER_114_600 ();
 FILLCELL_X2 FILLER_114_609 ();
 FILLCELL_X2 FILLER_114_632 ();
 FILLCELL_X8 FILLER_114_636 ();
 FILLCELL_X1 FILLER_114_644 ();
 FILLCELL_X4 FILLER_114_655 ();
 FILLCELL_X2 FILLER_114_659 ();
 FILLCELL_X1 FILLER_114_661 ();
 FILLCELL_X4 FILLER_114_689 ();
 FILLCELL_X2 FILLER_114_693 ();
 FILLCELL_X1 FILLER_114_695 ();
 FILLCELL_X2 FILLER_114_703 ();
 FILLCELL_X1 FILLER_114_710 ();
 FILLCELL_X4 FILLER_114_731 ();
 FILLCELL_X2 FILLER_114_735 ();
 FILLCELL_X1 FILLER_114_737 ();
 FILLCELL_X1 FILLER_114_758 ();
 FILLCELL_X2 FILLER_114_782 ();
 FILLCELL_X1 FILLER_114_784 ();
 FILLCELL_X2 FILLER_114_803 ();
 FILLCELL_X2 FILLER_114_823 ();
 FILLCELL_X1 FILLER_114_839 ();
 FILLCELL_X4 FILLER_114_865 ();
 FILLCELL_X1 FILLER_114_884 ();
 FILLCELL_X1 FILLER_114_889 ();
 FILLCELL_X2 FILLER_114_895 ();
 FILLCELL_X2 FILLER_114_908 ();
 FILLCELL_X4 FILLER_114_929 ();
 FILLCELL_X2 FILLER_114_933 ();
 FILLCELL_X2 FILLER_114_945 ();
 FILLCELL_X1 FILLER_114_947 ();
 FILLCELL_X4 FILLER_114_973 ();
 FILLCELL_X1 FILLER_114_977 ();
 FILLCELL_X8 FILLER_114_1000 ();
 FILLCELL_X1 FILLER_114_1008 ();
 FILLCELL_X4 FILLER_114_1031 ();
 FILLCELL_X4 FILLER_114_1057 ();
 FILLCELL_X1 FILLER_114_1061 ();
 FILLCELL_X1 FILLER_114_1065 ();
 FILLCELL_X16 FILLER_114_1081 ();
 FILLCELL_X1 FILLER_114_1097 ();
 FILLCELL_X8 FILLER_114_1100 ();
 FILLCELL_X4 FILLER_114_1108 ();
 FILLCELL_X8 FILLER_114_1133 ();
 FILLCELL_X4 FILLER_114_1141 ();
 FILLCELL_X2 FILLER_114_1145 ();
 FILLCELL_X4 FILLER_114_1178 ();
 FILLCELL_X2 FILLER_114_1213 ();
 FILLCELL_X1 FILLER_114_1215 ();
 FILLCELL_X8 FILLER_114_1221 ();
 FILLCELL_X4 FILLER_114_1229 ();
 FILLCELL_X2 FILLER_114_1233 ();
 FILLCELL_X1 FILLER_114_1235 ();
 FILLCELL_X4 FILLER_114_1239 ();
 FILLCELL_X2 FILLER_114_1243 ();
 FILLCELL_X1 FILLER_114_1245 ();
 FILLCELL_X16 FILLER_115_35 ();
 FILLCELL_X2 FILLER_115_51 ();
 FILLCELL_X1 FILLER_115_53 ();
 FILLCELL_X4 FILLER_115_74 ();
 FILLCELL_X16 FILLER_115_119 ();
 FILLCELL_X2 FILLER_115_135 ();
 FILLCELL_X8 FILLER_115_144 ();
 FILLCELL_X4 FILLER_115_152 ();
 FILLCELL_X2 FILLER_115_156 ();
 FILLCELL_X1 FILLER_115_158 ();
 FILLCELL_X4 FILLER_115_179 ();
 FILLCELL_X1 FILLER_115_209 ();
 FILLCELL_X2 FILLER_115_213 ();
 FILLCELL_X1 FILLER_115_215 ();
 FILLCELL_X4 FILLER_115_220 ();
 FILLCELL_X1 FILLER_115_224 ();
 FILLCELL_X2 FILLER_115_228 ();
 FILLCELL_X1 FILLER_115_230 ();
 FILLCELL_X4 FILLER_115_241 ();
 FILLCELL_X2 FILLER_115_245 ();
 FILLCELL_X1 FILLER_115_247 ();
 FILLCELL_X2 FILLER_115_252 ();
 FILLCELL_X1 FILLER_115_260 ();
 FILLCELL_X4 FILLER_115_276 ();
 FILLCELL_X1 FILLER_115_280 ();
 FILLCELL_X8 FILLER_115_301 ();
 FILLCELL_X2 FILLER_115_309 ();
 FILLCELL_X1 FILLER_115_311 ();
 FILLCELL_X4 FILLER_115_316 ();
 FILLCELL_X4 FILLER_115_323 ();
 FILLCELL_X2 FILLER_115_340 ();
 FILLCELL_X1 FILLER_115_354 ();
 FILLCELL_X4 FILLER_115_409 ();
 FILLCELL_X2 FILLER_115_413 ();
 FILLCELL_X2 FILLER_115_422 ();
 FILLCELL_X8 FILLER_115_435 ();
 FILLCELL_X2 FILLER_115_443 ();
 FILLCELL_X1 FILLER_115_445 ();
 FILLCELL_X2 FILLER_115_453 ();
 FILLCELL_X1 FILLER_115_455 ();
 FILLCELL_X4 FILLER_115_466 ();
 FILLCELL_X16 FILLER_115_530 ();
 FILLCELL_X4 FILLER_115_546 ();
 FILLCELL_X1 FILLER_115_550 ();
 FILLCELL_X8 FILLER_115_558 ();
 FILLCELL_X2 FILLER_115_578 ();
 FILLCELL_X1 FILLER_115_594 ();
 FILLCELL_X16 FILLER_115_615 ();
 FILLCELL_X8 FILLER_115_631 ();
 FILLCELL_X1 FILLER_115_662 ();
 FILLCELL_X4 FILLER_115_668 ();
 FILLCELL_X2 FILLER_115_672 ();
 FILLCELL_X8 FILLER_115_688 ();
 FILLCELL_X2 FILLER_115_696 ();
 FILLCELL_X1 FILLER_115_702 ();
 FILLCELL_X1 FILLER_115_712 ();
 FILLCELL_X8 FILLER_115_720 ();
 FILLCELL_X4 FILLER_115_728 ();
 FILLCELL_X2 FILLER_115_732 ();
 FILLCELL_X1 FILLER_115_746 ();
 FILLCELL_X4 FILLER_115_757 ();
 FILLCELL_X2 FILLER_115_761 ();
 FILLCELL_X2 FILLER_115_772 ();
 FILLCELL_X1 FILLER_115_774 ();
 FILLCELL_X2 FILLER_115_784 ();
 FILLCELL_X1 FILLER_115_786 ();
 FILLCELL_X1 FILLER_115_790 ();
 FILLCELL_X1 FILLER_115_798 ();
 FILLCELL_X1 FILLER_115_804 ();
 FILLCELL_X1 FILLER_115_809 ();
 FILLCELL_X2 FILLER_115_814 ();
 FILLCELL_X1 FILLER_115_834 ();
 FILLCELL_X2 FILLER_115_842 ();
 FILLCELL_X1 FILLER_115_844 ();
 FILLCELL_X2 FILLER_115_850 ();
 FILLCELL_X8 FILLER_115_866 ();
 FILLCELL_X4 FILLER_115_874 ();
 FILLCELL_X2 FILLER_115_878 ();
 FILLCELL_X1 FILLER_115_887 ();
 FILLCELL_X1 FILLER_115_897 ();
 FILLCELL_X4 FILLER_115_907 ();
 FILLCELL_X2 FILLER_115_964 ();
 FILLCELL_X1 FILLER_115_966 ();
 FILLCELL_X8 FILLER_115_971 ();
 FILLCELL_X4 FILLER_115_979 ();
 FILLCELL_X2 FILLER_115_987 ();
 FILLCELL_X1 FILLER_115_989 ();
 FILLCELL_X2 FILLER_115_1000 ();
 FILLCELL_X32 FILLER_115_1034 ();
 FILLCELL_X16 FILLER_115_1066 ();
 FILLCELL_X4 FILLER_115_1082 ();
 FILLCELL_X2 FILLER_115_1093 ();
 FILLCELL_X8 FILLER_115_1115 ();
 FILLCELL_X2 FILLER_115_1123 ();
 FILLCELL_X4 FILLER_115_1136 ();
 FILLCELL_X2 FILLER_115_1140 ();
 FILLCELL_X1 FILLER_115_1167 ();
 FILLCELL_X2 FILLER_115_1192 ();
 FILLCELL_X16 FILLER_115_1218 ();
 FILLCELL_X2 FILLER_115_1234 ();
 FILLCELL_X1 FILLER_115_1236 ();
 FILLCELL_X2 FILLER_115_1240 ();
 FILLCELL_X8 FILLER_115_1245 ();
 FILLCELL_X2 FILLER_115_1253 ();
 FILLCELL_X8 FILLER_116_21 ();
 FILLCELL_X4 FILLER_116_29 ();
 FILLCELL_X1 FILLER_116_60 ();
 FILLCELL_X4 FILLER_116_98 ();
 FILLCELL_X4 FILLER_116_109 ();
 FILLCELL_X2 FILLER_116_120 ();
 FILLCELL_X1 FILLER_116_122 ();
 FILLCELL_X4 FILLER_116_150 ();
 FILLCELL_X2 FILLER_116_154 ();
 FILLCELL_X8 FILLER_116_170 ();
 FILLCELL_X1 FILLER_116_178 ();
 FILLCELL_X1 FILLER_116_193 ();
 FILLCELL_X4 FILLER_116_208 ();
 FILLCELL_X2 FILLER_116_232 ();
 FILLCELL_X2 FILLER_116_238 ();
 FILLCELL_X16 FILLER_116_266 ();
 FILLCELL_X2 FILLER_116_282 ();
 FILLCELL_X1 FILLER_116_291 ();
 FILLCELL_X1 FILLER_116_295 ();
 FILLCELL_X16 FILLER_116_312 ();
 FILLCELL_X2 FILLER_116_328 ();
 FILLCELL_X1 FILLER_116_330 ();
 FILLCELL_X4 FILLER_116_351 ();
 FILLCELL_X16 FILLER_116_362 ();
 FILLCELL_X8 FILLER_116_378 ();
 FILLCELL_X1 FILLER_116_386 ();
 FILLCELL_X1 FILLER_116_392 ();
 FILLCELL_X1 FILLER_116_397 ();
 FILLCELL_X2 FILLER_116_405 ();
 FILLCELL_X2 FILLER_116_427 ();
 FILLCELL_X2 FILLER_116_436 ();
 FILLCELL_X1 FILLER_116_438 ();
 FILLCELL_X1 FILLER_116_453 ();
 FILLCELL_X1 FILLER_116_461 ();
 FILLCELL_X2 FILLER_116_469 ();
 FILLCELL_X1 FILLER_116_471 ();
 FILLCELL_X2 FILLER_116_485 ();
 FILLCELL_X1 FILLER_116_487 ();
 FILLCELL_X1 FILLER_116_495 ();
 FILLCELL_X8 FILLER_116_530 ();
 FILLCELL_X4 FILLER_116_538 ();
 FILLCELL_X2 FILLER_116_542 ();
 FILLCELL_X1 FILLER_116_544 ();
 FILLCELL_X32 FILLER_116_597 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X16 FILLER_116_632 ();
 FILLCELL_X2 FILLER_116_648 ();
 FILLCELL_X1 FILLER_116_650 ();
 FILLCELL_X1 FILLER_116_658 ();
 FILLCELL_X16 FILLER_116_699 ();
 FILLCELL_X8 FILLER_116_715 ();
 FILLCELL_X1 FILLER_116_723 ();
 FILLCELL_X4 FILLER_116_731 ();
 FILLCELL_X1 FILLER_116_735 ();
 FILLCELL_X1 FILLER_116_747 ();
 FILLCELL_X8 FILLER_116_768 ();
 FILLCELL_X1 FILLER_116_776 ();
 FILLCELL_X2 FILLER_116_782 ();
 FILLCELL_X4 FILLER_116_843 ();
 FILLCELL_X1 FILLER_116_854 ();
 FILLCELL_X2 FILLER_116_867 ();
 FILLCELL_X1 FILLER_116_869 ();
 FILLCELL_X1 FILLER_116_874 ();
 FILLCELL_X4 FILLER_116_892 ();
 FILLCELL_X4 FILLER_116_901 ();
 FILLCELL_X2 FILLER_116_905 ();
 FILLCELL_X1 FILLER_116_928 ();
 FILLCELL_X8 FILLER_116_941 ();
 FILLCELL_X2 FILLER_116_979 ();
 FILLCELL_X1 FILLER_116_985 ();
 FILLCELL_X1 FILLER_116_997 ();
 FILLCELL_X4 FILLER_116_1002 ();
 FILLCELL_X1 FILLER_116_1010 ();
 FILLCELL_X2 FILLER_116_1038 ();
 FILLCELL_X2 FILLER_116_1048 ();
 FILLCELL_X4 FILLER_116_1055 ();
 FILLCELL_X1 FILLER_116_1059 ();
 FILLCELL_X1 FILLER_116_1105 ();
 FILLCELL_X1 FILLER_116_1133 ();
 FILLCELL_X16 FILLER_116_1154 ();
 FILLCELL_X4 FILLER_116_1170 ();
 FILLCELL_X2 FILLER_116_1174 ();
 FILLCELL_X1 FILLER_116_1176 ();
 FILLCELL_X4 FILLER_116_1184 ();
 FILLCELL_X1 FILLER_116_1188 ();
 FILLCELL_X4 FILLER_116_1210 ();
 FILLCELL_X4 FILLER_116_1217 ();
 FILLCELL_X2 FILLER_116_1221 ();
 FILLCELL_X8 FILLER_116_1226 ();
 FILLCELL_X2 FILLER_116_1234 ();
 FILLCELL_X16 FILLER_116_1239 ();
 FILLCELL_X8 FILLER_117_1 ();
 FILLCELL_X2 FILLER_117_9 ();
 FILLCELL_X1 FILLER_117_18 ();
 FILLCELL_X4 FILLER_117_39 ();
 FILLCELL_X2 FILLER_117_76 ();
 FILLCELL_X16 FILLER_117_92 ();
 FILLCELL_X2 FILLER_117_108 ();
 FILLCELL_X1 FILLER_117_110 ();
 FILLCELL_X2 FILLER_117_118 ();
 FILLCELL_X4 FILLER_117_127 ();
 FILLCELL_X2 FILLER_117_131 ();
 FILLCELL_X1 FILLER_117_133 ();
 FILLCELL_X4 FILLER_117_148 ();
 FILLCELL_X2 FILLER_117_152 ();
 FILLCELL_X1 FILLER_117_154 ();
 FILLCELL_X4 FILLER_117_203 ();
 FILLCELL_X2 FILLER_117_207 ();
 FILLCELL_X8 FILLER_117_223 ();
 FILLCELL_X2 FILLER_117_231 ();
 FILLCELL_X1 FILLER_117_233 ();
 FILLCELL_X8 FILLER_117_241 ();
 FILLCELL_X1 FILLER_117_249 ();
 FILLCELL_X2 FILLER_117_253 ();
 FILLCELL_X1 FILLER_117_255 ();
 FILLCELL_X2 FILLER_117_301 ();
 FILLCELL_X4 FILLER_117_314 ();
 FILLCELL_X1 FILLER_117_318 ();
 FILLCELL_X2 FILLER_117_323 ();
 FILLCELL_X4 FILLER_117_330 ();
 FILLCELL_X2 FILLER_117_334 ();
 FILLCELL_X1 FILLER_117_343 ();
 FILLCELL_X1 FILLER_117_364 ();
 FILLCELL_X1 FILLER_117_375 ();
 FILLCELL_X1 FILLER_117_382 ();
 FILLCELL_X4 FILLER_117_433 ();
 FILLCELL_X2 FILLER_117_444 ();
 FILLCELL_X2 FILLER_117_453 ();
 FILLCELL_X1 FILLER_117_455 ();
 FILLCELL_X4 FILLER_117_525 ();
 FILLCELL_X1 FILLER_117_529 ();
 FILLCELL_X2 FILLER_117_551 ();
 FILLCELL_X4 FILLER_117_560 ();
 FILLCELL_X1 FILLER_117_564 ();
 FILLCELL_X8 FILLER_117_586 ();
 FILLCELL_X1 FILLER_117_594 ();
 FILLCELL_X2 FILLER_117_622 ();
 FILLCELL_X4 FILLER_117_643 ();
 FILLCELL_X1 FILLER_117_647 ();
 FILLCELL_X2 FILLER_117_655 ();
 FILLCELL_X1 FILLER_117_664 ();
 FILLCELL_X2 FILLER_117_672 ();
 FILLCELL_X8 FILLER_117_681 ();
 FILLCELL_X4 FILLER_117_689 ();
 FILLCELL_X2 FILLER_117_693 ();
 FILLCELL_X8 FILLER_117_723 ();
 FILLCELL_X4 FILLER_117_742 ();
 FILLCELL_X1 FILLER_117_746 ();
 FILLCELL_X8 FILLER_117_754 ();
 FILLCELL_X4 FILLER_117_762 ();
 FILLCELL_X1 FILLER_117_771 ();
 FILLCELL_X8 FILLER_117_779 ();
 FILLCELL_X1 FILLER_117_787 ();
 FILLCELL_X8 FILLER_117_793 ();
 FILLCELL_X4 FILLER_117_801 ();
 FILLCELL_X2 FILLER_117_805 ();
 FILLCELL_X1 FILLER_117_807 ();
 FILLCELL_X2 FILLER_117_824 ();
 FILLCELL_X4 FILLER_117_830 ();
 FILLCELL_X2 FILLER_117_842 ();
 FILLCELL_X1 FILLER_117_844 ();
 FILLCELL_X4 FILLER_117_856 ();
 FILLCELL_X1 FILLER_117_860 ();
 FILLCELL_X2 FILLER_117_874 ();
 FILLCELL_X1 FILLER_117_876 ();
 FILLCELL_X4 FILLER_117_921 ();
 FILLCELL_X8 FILLER_117_928 ();
 FILLCELL_X4 FILLER_117_936 ();
 FILLCELL_X2 FILLER_117_961 ();
 FILLCELL_X4 FILLER_117_973 ();
 FILLCELL_X2 FILLER_117_977 ();
 FILLCELL_X4 FILLER_117_985 ();
 FILLCELL_X2 FILLER_117_992 ();
 FILLCELL_X1 FILLER_117_994 ();
 FILLCELL_X8 FILLER_117_1005 ();
 FILLCELL_X4 FILLER_117_1013 ();
 FILLCELL_X2 FILLER_117_1017 ();
 FILLCELL_X2 FILLER_117_1033 ();
 FILLCELL_X1 FILLER_117_1042 ();
 FILLCELL_X4 FILLER_117_1052 ();
 FILLCELL_X2 FILLER_117_1056 ();
 FILLCELL_X8 FILLER_117_1075 ();
 FILLCELL_X2 FILLER_117_1083 ();
 FILLCELL_X1 FILLER_117_1085 ();
 FILLCELL_X16 FILLER_117_1108 ();
 FILLCELL_X4 FILLER_117_1124 ();
 FILLCELL_X8 FILLER_117_1133 ();
 FILLCELL_X1 FILLER_117_1141 ();
 FILLCELL_X4 FILLER_117_1173 ();
 FILLCELL_X1 FILLER_117_1177 ();
 FILLCELL_X4 FILLER_117_1185 ();
 FILLCELL_X4 FILLER_117_1196 ();
 FILLCELL_X2 FILLER_117_1200 ();
 FILLCELL_X1 FILLER_117_1202 ();
 FILLCELL_X4 FILLER_117_1220 ();
 FILLCELL_X1 FILLER_117_1224 ();
 FILLCELL_X2 FILLER_117_1228 ();
 FILLCELL_X1 FILLER_117_1230 ();
 FILLCELL_X16 FILLER_117_1234 ();
 FILLCELL_X4 FILLER_117_1250 ();
 FILLCELL_X1 FILLER_117_1254 ();
 FILLCELL_X16 FILLER_118_1 ();
 FILLCELL_X1 FILLER_118_17 ();
 FILLCELL_X2 FILLER_118_38 ();
 FILLCELL_X4 FILLER_118_59 ();
 FILLCELL_X1 FILLER_118_63 ();
 FILLCELL_X2 FILLER_118_71 ();
 FILLCELL_X2 FILLER_118_87 ();
 FILLCELL_X4 FILLER_118_143 ();
 FILLCELL_X1 FILLER_118_147 ();
 FILLCELL_X8 FILLER_118_168 ();
 FILLCELL_X1 FILLER_118_194 ();
 FILLCELL_X2 FILLER_118_199 ();
 FILLCELL_X1 FILLER_118_201 ();
 FILLCELL_X8 FILLER_118_228 ();
 FILLCELL_X4 FILLER_118_236 ();
 FILLCELL_X2 FILLER_118_244 ();
 FILLCELL_X8 FILLER_118_249 ();
 FILLCELL_X2 FILLER_118_257 ();
 FILLCELL_X8 FILLER_118_272 ();
 FILLCELL_X2 FILLER_118_280 ();
 FILLCELL_X1 FILLER_118_282 ();
 FILLCELL_X2 FILLER_118_287 ();
 FILLCELL_X1 FILLER_118_289 ();
 FILLCELL_X2 FILLER_118_293 ();
 FILLCELL_X1 FILLER_118_302 ();
 FILLCELL_X4 FILLER_118_313 ();
 FILLCELL_X1 FILLER_118_317 ();
 FILLCELL_X16 FILLER_118_338 ();
 FILLCELL_X4 FILLER_118_354 ();
 FILLCELL_X4 FILLER_118_365 ();
 FILLCELL_X1 FILLER_118_369 ();
 FILLCELL_X16 FILLER_118_385 ();
 FILLCELL_X8 FILLER_118_401 ();
 FILLCELL_X4 FILLER_118_409 ();
 FILLCELL_X2 FILLER_118_413 ();
 FILLCELL_X1 FILLER_118_415 ();
 FILLCELL_X4 FILLER_118_431 ();
 FILLCELL_X1 FILLER_118_435 ();
 FILLCELL_X4 FILLER_118_446 ();
 FILLCELL_X1 FILLER_118_450 ();
 FILLCELL_X2 FILLER_118_470 ();
 FILLCELL_X1 FILLER_118_472 ();
 FILLCELL_X2 FILLER_118_486 ();
 FILLCELL_X1 FILLER_118_488 ();
 FILLCELL_X4 FILLER_118_498 ();
 FILLCELL_X2 FILLER_118_502 ();
 FILLCELL_X1 FILLER_118_504 ();
 FILLCELL_X1 FILLER_118_537 ();
 FILLCELL_X8 FILLER_118_571 ();
 FILLCELL_X2 FILLER_118_579 ();
 FILLCELL_X4 FILLER_118_588 ();
 FILLCELL_X2 FILLER_118_599 ();
 FILLCELL_X8 FILLER_118_621 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X2 FILLER_118_632 ();
 FILLCELL_X1 FILLER_118_634 ();
 FILLCELL_X8 FILLER_118_639 ();
 FILLCELL_X1 FILLER_118_647 ();
 FILLCELL_X4 FILLER_118_720 ();
 FILLCELL_X1 FILLER_118_724 ();
 FILLCELL_X4 FILLER_118_747 ();
 FILLCELL_X4 FILLER_118_758 ();
 FILLCELL_X4 FILLER_118_803 ();
 FILLCELL_X2 FILLER_118_807 ();
 FILLCELL_X2 FILLER_118_826 ();
 FILLCELL_X4 FILLER_118_833 ();
 FILLCELL_X1 FILLER_118_868 ();
 FILLCELL_X1 FILLER_118_880 ();
 FILLCELL_X1 FILLER_118_894 ();
 FILLCELL_X1 FILLER_118_897 ();
 FILLCELL_X1 FILLER_118_910 ();
 FILLCELL_X2 FILLER_118_920 ();
 FILLCELL_X4 FILLER_118_929 ();
 FILLCELL_X2 FILLER_118_933 ();
 FILLCELL_X4 FILLER_118_939 ();
 FILLCELL_X2 FILLER_118_943 ();
 FILLCELL_X8 FILLER_118_955 ();
 FILLCELL_X4 FILLER_118_963 ();
 FILLCELL_X2 FILLER_118_971 ();
 FILLCELL_X8 FILLER_118_990 ();
 FILLCELL_X1 FILLER_118_998 ();
 FILLCELL_X1 FILLER_118_1029 ();
 FILLCELL_X32 FILLER_118_1033 ();
 FILLCELL_X4 FILLER_118_1065 ();
 FILLCELL_X1 FILLER_118_1100 ();
 FILLCELL_X2 FILLER_118_1108 ();
 FILLCELL_X2 FILLER_118_1114 ();
 FILLCELL_X1 FILLER_118_1116 ();
 FILLCELL_X4 FILLER_118_1141 ();
 FILLCELL_X2 FILLER_118_1145 ();
 FILLCELL_X1 FILLER_118_1147 ();
 FILLCELL_X8 FILLER_118_1153 ();
 FILLCELL_X2 FILLER_118_1161 ();
 FILLCELL_X1 FILLER_118_1163 ();
 FILLCELL_X2 FILLER_118_1171 ();
 FILLCELL_X1 FILLER_118_1173 ();
 FILLCELL_X16 FILLER_118_1208 ();
 FILLCELL_X2 FILLER_118_1224 ();
 FILLCELL_X1 FILLER_118_1226 ();
 FILLCELL_X8 FILLER_118_1233 ();
 FILLCELL_X8 FILLER_118_1244 ();
 FILLCELL_X2 FILLER_118_1252 ();
 FILLCELL_X1 FILLER_118_1254 ();
 FILLCELL_X8 FILLER_119_1 ();
 FILLCELL_X4 FILLER_119_9 ();
 FILLCELL_X1 FILLER_119_13 ();
 FILLCELL_X4 FILLER_119_21 ();
 FILLCELL_X2 FILLER_119_67 ();
 FILLCELL_X8 FILLER_119_90 ();
 FILLCELL_X2 FILLER_119_98 ();
 FILLCELL_X1 FILLER_119_100 ();
 FILLCELL_X8 FILLER_119_108 ();
 FILLCELL_X2 FILLER_119_116 ();
 FILLCELL_X1 FILLER_119_118 ();
 FILLCELL_X8 FILLER_119_126 ();
 FILLCELL_X2 FILLER_119_134 ();
 FILLCELL_X4 FILLER_119_143 ();
 FILLCELL_X1 FILLER_119_147 ();
 FILLCELL_X2 FILLER_119_155 ();
 FILLCELL_X1 FILLER_119_255 ();
 FILLCELL_X1 FILLER_119_263 ();
 FILLCELL_X1 FILLER_119_268 ();
 FILLCELL_X1 FILLER_119_293 ();
 FILLCELL_X1 FILLER_119_301 ();
 FILLCELL_X4 FILLER_119_313 ();
 FILLCELL_X1 FILLER_119_317 ();
 FILLCELL_X32 FILLER_119_325 ();
 FILLCELL_X4 FILLER_119_377 ();
 FILLCELL_X2 FILLER_119_395 ();
 FILLCELL_X1 FILLER_119_397 ();
 FILLCELL_X2 FILLER_119_425 ();
 FILLCELL_X2 FILLER_119_434 ();
 FILLCELL_X1 FILLER_119_436 ();
 FILLCELL_X1 FILLER_119_444 ();
 FILLCELL_X2 FILLER_119_466 ();
 FILLCELL_X1 FILLER_119_468 ();
 FILLCELL_X1 FILLER_119_472 ();
 FILLCELL_X1 FILLER_119_480 ();
 FILLCELL_X4 FILLER_119_485 ();
 FILLCELL_X1 FILLER_119_489 ();
 FILLCELL_X2 FILLER_119_526 ();
 FILLCELL_X1 FILLER_119_528 ();
 FILLCELL_X32 FILLER_119_542 ();
 FILLCELL_X2 FILLER_119_574 ();
 FILLCELL_X1 FILLER_119_576 ();
 FILLCELL_X4 FILLER_119_660 ();
 FILLCELL_X1 FILLER_119_664 ();
 FILLCELL_X2 FILLER_119_672 ();
 FILLCELL_X8 FILLER_119_681 ();
 FILLCELL_X4 FILLER_119_689 ();
 FILLCELL_X1 FILLER_119_693 ();
 FILLCELL_X4 FILLER_119_708 ();
 FILLCELL_X2 FILLER_119_712 ();
 FILLCELL_X1 FILLER_119_714 ();
 FILLCELL_X1 FILLER_119_722 ();
 FILLCELL_X1 FILLER_119_730 ();
 FILLCELL_X1 FILLER_119_738 ();
 FILLCELL_X1 FILLER_119_746 ();
 FILLCELL_X16 FILLER_119_767 ();
 FILLCELL_X2 FILLER_119_783 ();
 FILLCELL_X1 FILLER_119_785 ();
 FILLCELL_X2 FILLER_119_816 ();
 FILLCELL_X8 FILLER_119_825 ();
 FILLCELL_X1 FILLER_119_833 ();
 FILLCELL_X4 FILLER_119_843 ();
 FILLCELL_X2 FILLER_119_847 ();
 FILLCELL_X1 FILLER_119_849 ();
 FILLCELL_X8 FILLER_119_857 ();
 FILLCELL_X8 FILLER_119_872 ();
 FILLCELL_X2 FILLER_119_880 ();
 FILLCELL_X2 FILLER_119_904 ();
 FILLCELL_X1 FILLER_119_906 ();
 FILLCELL_X1 FILLER_119_955 ();
 FILLCELL_X1 FILLER_119_967 ();
 FILLCELL_X2 FILLER_119_971 ();
 FILLCELL_X8 FILLER_119_976 ();
 FILLCELL_X4 FILLER_119_984 ();
 FILLCELL_X8 FILLER_119_991 ();
 FILLCELL_X2 FILLER_119_999 ();
 FILLCELL_X16 FILLER_119_1004 ();
 FILLCELL_X8 FILLER_119_1020 ();
 FILLCELL_X2 FILLER_119_1031 ();
 FILLCELL_X1 FILLER_119_1033 ();
 FILLCELL_X8 FILLER_119_1057 ();
 FILLCELL_X1 FILLER_119_1065 ();
 FILLCELL_X4 FILLER_119_1069 ();
 FILLCELL_X2 FILLER_119_1080 ();
 FILLCELL_X4 FILLER_119_1098 ();
 FILLCELL_X2 FILLER_119_1102 ();
 FILLCELL_X1 FILLER_119_1104 ();
 FILLCELL_X8 FILLER_119_1112 ();
 FILLCELL_X1 FILLER_119_1120 ();
 FILLCELL_X2 FILLER_119_1123 ();
 FILLCELL_X4 FILLER_119_1155 ();
 FILLCELL_X1 FILLER_119_1159 ();
 FILLCELL_X32 FILLER_119_1180 ();
 FILLCELL_X16 FILLER_119_1212 ();
 FILLCELL_X8 FILLER_119_1228 ();
 FILLCELL_X1 FILLER_119_1236 ();
 FILLCELL_X8 FILLER_119_1240 ();
 FILLCELL_X4 FILLER_119_1248 ();
 FILLCELL_X2 FILLER_119_1252 ();
 FILLCELL_X1 FILLER_119_1254 ();
 FILLCELL_X4 FILLER_120_1 ();
 FILLCELL_X2 FILLER_120_5 ();
 FILLCELL_X1 FILLER_120_7 ();
 FILLCELL_X1 FILLER_120_15 ();
 FILLCELL_X16 FILLER_120_43 ();
 FILLCELL_X4 FILLER_120_86 ();
 FILLCELL_X2 FILLER_120_90 ();
 FILLCELL_X2 FILLER_120_150 ();
 FILLCELL_X2 FILLER_120_172 ();
 FILLCELL_X16 FILLER_120_176 ();
 FILLCELL_X1 FILLER_120_192 ();
 FILLCELL_X2 FILLER_120_202 ();
 FILLCELL_X1 FILLER_120_204 ();
 FILLCELL_X16 FILLER_120_222 ();
 FILLCELL_X8 FILLER_120_238 ();
 FILLCELL_X1 FILLER_120_246 ();
 FILLCELL_X2 FILLER_120_261 ();
 FILLCELL_X16 FILLER_120_270 ();
 FILLCELL_X1 FILLER_120_286 ();
 FILLCELL_X1 FILLER_120_291 ();
 FILLCELL_X4 FILLER_120_299 ();
 FILLCELL_X1 FILLER_120_303 ();
 FILLCELL_X2 FILLER_120_314 ();
 FILLCELL_X2 FILLER_120_336 ();
 FILLCELL_X1 FILLER_120_338 ();
 FILLCELL_X1 FILLER_120_366 ();
 FILLCELL_X2 FILLER_120_380 ();
 FILLCELL_X1 FILLER_120_386 ();
 FILLCELL_X4 FILLER_120_393 ();
 FILLCELL_X2 FILLER_120_397 ();
 FILLCELL_X4 FILLER_120_441 ();
 FILLCELL_X8 FILLER_120_512 ();
 FILLCELL_X1 FILLER_120_520 ();
 FILLCELL_X2 FILLER_120_541 ();
 FILLCELL_X4 FILLER_120_550 ();
 FILLCELL_X2 FILLER_120_554 ();
 FILLCELL_X4 FILLER_120_563 ();
 FILLCELL_X2 FILLER_120_567 ();
 FILLCELL_X2 FILLER_120_594 ();
 FILLCELL_X2 FILLER_120_603 ();
 FILLCELL_X1 FILLER_120_630 ();
 FILLCELL_X2 FILLER_120_632 ();
 FILLCELL_X8 FILLER_120_638 ();
 FILLCELL_X4 FILLER_120_646 ();
 FILLCELL_X4 FILLER_120_670 ();
 FILLCELL_X2 FILLER_120_674 ();
 FILLCELL_X1 FILLER_120_703 ();
 FILLCELL_X8 FILLER_120_731 ();
 FILLCELL_X2 FILLER_120_739 ();
 FILLCELL_X1 FILLER_120_761 ();
 FILLCELL_X4 FILLER_120_804 ();
 FILLCELL_X2 FILLER_120_808 ();
 FILLCELL_X4 FILLER_120_831 ();
 FILLCELL_X2 FILLER_120_835 ();
 FILLCELL_X4 FILLER_120_862 ();
 FILLCELL_X2 FILLER_120_866 ();
 FILLCELL_X4 FILLER_120_875 ();
 FILLCELL_X1 FILLER_120_879 ();
 FILLCELL_X2 FILLER_120_883 ();
 FILLCELL_X1 FILLER_120_889 ();
 FILLCELL_X8 FILLER_120_897 ();
 FILLCELL_X1 FILLER_120_905 ();
 FILLCELL_X2 FILLER_120_912 ();
 FILLCELL_X1 FILLER_120_914 ();
 FILLCELL_X1 FILLER_120_924 ();
 FILLCELL_X4 FILLER_120_929 ();
 FILLCELL_X1 FILLER_120_933 ();
 FILLCELL_X4 FILLER_120_947 ();
 FILLCELL_X4 FILLER_120_955 ();
 FILLCELL_X2 FILLER_120_973 ();
 FILLCELL_X1 FILLER_120_975 ();
 FILLCELL_X1 FILLER_120_985 ();
 FILLCELL_X4 FILLER_120_996 ();
 FILLCELL_X2 FILLER_120_1000 ();
 FILLCELL_X4 FILLER_120_1007 ();
 FILLCELL_X2 FILLER_120_1021 ();
 FILLCELL_X1 FILLER_120_1032 ();
 FILLCELL_X8 FILLER_120_1040 ();
 FILLCELL_X1 FILLER_120_1048 ();
 FILLCELL_X2 FILLER_120_1072 ();
 FILLCELL_X1 FILLER_120_1098 ();
 FILLCELL_X2 FILLER_120_1123 ();
 FILLCELL_X1 FILLER_120_1125 ();
 FILLCELL_X4 FILLER_120_1130 ();
 FILLCELL_X2 FILLER_120_1134 ();
 FILLCELL_X8 FILLER_120_1162 ();
 FILLCELL_X1 FILLER_120_1170 ();
 FILLCELL_X32 FILLER_120_1175 ();
 FILLCELL_X16 FILLER_120_1207 ();
 FILLCELL_X4 FILLER_120_1223 ();
 FILLCELL_X1 FILLER_120_1227 ();
 FILLCELL_X16 FILLER_120_1234 ();
 FILLCELL_X2 FILLER_120_1253 ();
 FILLCELL_X16 FILLER_121_1 ();
 FILLCELL_X8 FILLER_121_17 ();
 FILLCELL_X1 FILLER_121_25 ();
 FILLCELL_X16 FILLER_121_46 ();
 FILLCELL_X2 FILLER_121_69 ();
 FILLCELL_X1 FILLER_121_98 ();
 FILLCELL_X1 FILLER_121_113 ();
 FILLCELL_X2 FILLER_121_133 ();
 FILLCELL_X2 FILLER_121_138 ();
 FILLCELL_X2 FILLER_121_144 ();
 FILLCELL_X1 FILLER_121_146 ();
 FILLCELL_X1 FILLER_121_151 ();
 FILLCELL_X2 FILLER_121_159 ();
 FILLCELL_X1 FILLER_121_161 ();
 FILLCELL_X8 FILLER_121_210 ();
 FILLCELL_X2 FILLER_121_218 ();
 FILLCELL_X1 FILLER_121_220 ();
 FILLCELL_X1 FILLER_121_228 ();
 FILLCELL_X4 FILLER_121_243 ();
 FILLCELL_X4 FILLER_121_250 ();
 FILLCELL_X16 FILLER_121_261 ();
 FILLCELL_X1 FILLER_121_300 ();
 FILLCELL_X4 FILLER_121_326 ();
 FILLCELL_X2 FILLER_121_330 ();
 FILLCELL_X1 FILLER_121_332 ();
 FILLCELL_X2 FILLER_121_360 ();
 FILLCELL_X1 FILLER_121_362 ();
 FILLCELL_X1 FILLER_121_384 ();
 FILLCELL_X4 FILLER_121_399 ();
 FILLCELL_X2 FILLER_121_403 ();
 FILLCELL_X1 FILLER_121_405 ();
 FILLCELL_X2 FILLER_121_413 ();
 FILLCELL_X1 FILLER_121_415 ();
 FILLCELL_X8 FILLER_121_480 ();
 FILLCELL_X4 FILLER_121_502 ();
 FILLCELL_X2 FILLER_121_506 ();
 FILLCELL_X2 FILLER_121_513 ();
 FILLCELL_X4 FILLER_121_522 ();
 FILLCELL_X1 FILLER_121_526 ();
 FILLCELL_X4 FILLER_121_547 ();
 FILLCELL_X1 FILLER_121_551 ();
 FILLCELL_X4 FILLER_121_572 ();
 FILLCELL_X1 FILLER_121_583 ();
 FILLCELL_X4 FILLER_121_598 ();
 FILLCELL_X8 FILLER_121_609 ();
 FILLCELL_X2 FILLER_121_619 ();
 FILLCELL_X1 FILLER_121_621 ();
 FILLCELL_X4 FILLER_121_626 ();
 FILLCELL_X8 FILLER_121_640 ();
 FILLCELL_X1 FILLER_121_648 ();
 FILLCELL_X8 FILLER_121_656 ();
 FILLCELL_X4 FILLER_121_664 ();
 FILLCELL_X1 FILLER_121_668 ();
 FILLCELL_X4 FILLER_121_690 ();
 FILLCELL_X1 FILLER_121_694 ();
 FILLCELL_X8 FILLER_121_702 ();
 FILLCELL_X1 FILLER_121_710 ();
 FILLCELL_X16 FILLER_121_718 ();
 FILLCELL_X1 FILLER_121_734 ();
 FILLCELL_X8 FILLER_121_742 ();
 FILLCELL_X4 FILLER_121_750 ();
 FILLCELL_X4 FILLER_121_761 ();
 FILLCELL_X2 FILLER_121_765 ();
 FILLCELL_X1 FILLER_121_767 ();
 FILLCELL_X8 FILLER_121_775 ();
 FILLCELL_X4 FILLER_121_783 ();
 FILLCELL_X1 FILLER_121_787 ();
 FILLCELL_X2 FILLER_121_795 ();
 FILLCELL_X1 FILLER_121_797 ();
 FILLCELL_X8 FILLER_121_805 ();
 FILLCELL_X1 FILLER_121_813 ();
 FILLCELL_X4 FILLER_121_844 ();
 FILLCELL_X1 FILLER_121_848 ();
 FILLCELL_X2 FILLER_121_865 ();
 FILLCELL_X1 FILLER_121_867 ();
 FILLCELL_X2 FILLER_121_894 ();
 FILLCELL_X1 FILLER_121_896 ();
 FILLCELL_X1 FILLER_121_923 ();
 FILLCELL_X2 FILLER_121_944 ();
 FILLCELL_X1 FILLER_121_961 ();
 FILLCELL_X1 FILLER_121_965 ();
 FILLCELL_X1 FILLER_121_970 ();
 FILLCELL_X1 FILLER_121_974 ();
 FILLCELL_X1 FILLER_121_978 ();
 FILLCELL_X1 FILLER_121_990 ();
 FILLCELL_X1 FILLER_121_1013 ();
 FILLCELL_X1 FILLER_121_1018 ();
 FILLCELL_X1 FILLER_121_1023 ();
 FILLCELL_X2 FILLER_121_1042 ();
 FILLCELL_X1 FILLER_121_1049 ();
 FILLCELL_X2 FILLER_121_1054 ();
 FILLCELL_X8 FILLER_121_1071 ();
 FILLCELL_X2 FILLER_121_1079 ();
 FILLCELL_X1 FILLER_121_1084 ();
 FILLCELL_X1 FILLER_121_1094 ();
 FILLCELL_X4 FILLER_121_1097 ();
 FILLCELL_X2 FILLER_121_1101 ();
 FILLCELL_X1 FILLER_121_1103 ();
 FILLCELL_X2 FILLER_121_1108 ();
 FILLCELL_X2 FILLER_121_1141 ();
 FILLCELL_X32 FILLER_121_1179 ();
 FILLCELL_X16 FILLER_121_1211 ();
 FILLCELL_X4 FILLER_121_1227 ();
 FILLCELL_X8 FILLER_121_1234 ();
 FILLCELL_X1 FILLER_121_1245 ();
 FILLCELL_X4 FILLER_121_1249 ();
 FILLCELL_X2 FILLER_121_1253 ();
 FILLCELL_X16 FILLER_122_1 ();
 FILLCELL_X4 FILLER_122_17 ();
 FILLCELL_X1 FILLER_122_21 ();
 FILLCELL_X4 FILLER_122_29 ();
 FILLCELL_X2 FILLER_122_33 ();
 FILLCELL_X1 FILLER_122_35 ();
 FILLCELL_X16 FILLER_122_57 ();
 FILLCELL_X8 FILLER_122_73 ();
 FILLCELL_X1 FILLER_122_81 ();
 FILLCELL_X2 FILLER_122_116 ();
 FILLCELL_X8 FILLER_122_145 ();
 FILLCELL_X4 FILLER_122_153 ();
 FILLCELL_X2 FILLER_122_180 ();
 FILLCELL_X8 FILLER_122_186 ();
 FILLCELL_X2 FILLER_122_194 ();
 FILLCELL_X1 FILLER_122_196 ();
 FILLCELL_X2 FILLER_122_230 ();
 FILLCELL_X1 FILLER_122_252 ();
 FILLCELL_X2 FILLER_122_276 ();
 FILLCELL_X1 FILLER_122_278 ();
 FILLCELL_X16 FILLER_122_292 ();
 FILLCELL_X1 FILLER_122_308 ();
 FILLCELL_X2 FILLER_122_319 ();
 FILLCELL_X1 FILLER_122_321 ();
 FILLCELL_X4 FILLER_122_349 ();
 FILLCELL_X2 FILLER_122_353 ();
 FILLCELL_X1 FILLER_122_355 ();
 FILLCELL_X4 FILLER_122_376 ();
 FILLCELL_X4 FILLER_122_403 ();
 FILLCELL_X1 FILLER_122_407 ();
 FILLCELL_X8 FILLER_122_428 ();
 FILLCELL_X4 FILLER_122_443 ();
 FILLCELL_X1 FILLER_122_447 ();
 FILLCELL_X2 FILLER_122_455 ();
 FILLCELL_X2 FILLER_122_464 ();
 FILLCELL_X8 FILLER_122_504 ();
 FILLCELL_X4 FILLER_122_512 ();
 FILLCELL_X2 FILLER_122_516 ();
 FILLCELL_X2 FILLER_122_538 ();
 FILLCELL_X1 FILLER_122_540 ();
 FILLCELL_X16 FILLER_122_548 ();
 FILLCELL_X4 FILLER_122_564 ();
 FILLCELL_X1 FILLER_122_568 ();
 FILLCELL_X8 FILLER_122_576 ();
 FILLCELL_X1 FILLER_122_584 ();
 FILLCELL_X4 FILLER_122_590 ();
 FILLCELL_X2 FILLER_122_594 ();
 FILLCELL_X4 FILLER_122_616 ();
 FILLCELL_X2 FILLER_122_620 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X8 FILLER_122_639 ();
 FILLCELL_X1 FILLER_122_647 ();
 FILLCELL_X8 FILLER_122_668 ();
 FILLCELL_X2 FILLER_122_676 ();
 FILLCELL_X1 FILLER_122_689 ();
 FILLCELL_X4 FILLER_122_703 ();
 FILLCELL_X1 FILLER_122_707 ();
 FILLCELL_X4 FILLER_122_729 ();
 FILLCELL_X2 FILLER_122_733 ();
 FILLCELL_X1 FILLER_122_735 ();
 FILLCELL_X4 FILLER_122_756 ();
 FILLCELL_X4 FILLER_122_767 ();
 FILLCELL_X2 FILLER_122_771 ();
 FILLCELL_X1 FILLER_122_773 ();
 FILLCELL_X4 FILLER_122_779 ();
 FILLCELL_X1 FILLER_122_783 ();
 FILLCELL_X1 FILLER_122_798 ();
 FILLCELL_X2 FILLER_122_819 ();
 FILLCELL_X1 FILLER_122_821 ();
 FILLCELL_X16 FILLER_122_824 ();
 FILLCELL_X8 FILLER_122_840 ();
 FILLCELL_X1 FILLER_122_848 ();
 FILLCELL_X2 FILLER_122_853 ();
 FILLCELL_X2 FILLER_122_869 ();
 FILLCELL_X1 FILLER_122_871 ();
 FILLCELL_X2 FILLER_122_879 ();
 FILLCELL_X1 FILLER_122_881 ();
 FILLCELL_X2 FILLER_122_888 ();
 FILLCELL_X1 FILLER_122_894 ();
 FILLCELL_X1 FILLER_122_898 ();
 FILLCELL_X4 FILLER_122_907 ();
 FILLCELL_X4 FILLER_122_915 ();
 FILLCELL_X8 FILLER_122_926 ();
 FILLCELL_X8 FILLER_122_938 ();
 FILLCELL_X2 FILLER_122_946 ();
 FILLCELL_X1 FILLER_122_948 ();
 FILLCELL_X2 FILLER_122_952 ();
 FILLCELL_X1 FILLER_122_972 ();
 FILLCELL_X2 FILLER_122_987 ();
 FILLCELL_X1 FILLER_122_989 ();
 FILLCELL_X8 FILLER_122_1003 ();
 FILLCELL_X4 FILLER_122_1011 ();
 FILLCELL_X1 FILLER_122_1022 ();
 FILLCELL_X4 FILLER_122_1027 ();
 FILLCELL_X1 FILLER_122_1031 ();
 FILLCELL_X2 FILLER_122_1069 ();
 FILLCELL_X1 FILLER_122_1071 ();
 FILLCELL_X8 FILLER_122_1084 ();
 FILLCELL_X4 FILLER_122_1092 ();
 FILLCELL_X2 FILLER_122_1096 ();
 FILLCELL_X8 FILLER_122_1118 ();
 FILLCELL_X2 FILLER_122_1126 ();
 FILLCELL_X1 FILLER_122_1128 ();
 FILLCELL_X4 FILLER_122_1134 ();
 FILLCELL_X2 FILLER_122_1138 ();
 FILLCELL_X1 FILLER_122_1140 ();
 FILLCELL_X16 FILLER_122_1194 ();
 FILLCELL_X8 FILLER_122_1210 ();
 FILLCELL_X2 FILLER_122_1218 ();
 FILLCELL_X1 FILLER_122_1220 ();
 FILLCELL_X1 FILLER_122_1224 ();
 FILLCELL_X2 FILLER_122_1228 ();
 FILLCELL_X1 FILLER_122_1230 ();
 FILLCELL_X16 FILLER_122_1234 ();
 FILLCELL_X4 FILLER_122_1250 ();
 FILLCELL_X1 FILLER_122_1254 ();
 FILLCELL_X4 FILLER_123_1 ();
 FILLCELL_X2 FILLER_123_5 ();
 FILLCELL_X1 FILLER_123_7 ();
 FILLCELL_X2 FILLER_123_15 ();
 FILLCELL_X1 FILLER_123_17 ();
 FILLCELL_X4 FILLER_123_38 ();
 FILLCELL_X16 FILLER_123_49 ();
 FILLCELL_X8 FILLER_123_65 ();
 FILLCELL_X4 FILLER_123_73 ();
 FILLCELL_X16 FILLER_123_97 ();
 FILLCELL_X4 FILLER_123_113 ();
 FILLCELL_X4 FILLER_123_124 ();
 FILLCELL_X2 FILLER_123_128 ();
 FILLCELL_X4 FILLER_123_171 ();
 FILLCELL_X2 FILLER_123_193 ();
 FILLCELL_X4 FILLER_123_222 ();
 FILLCELL_X1 FILLER_123_226 ();
 FILLCELL_X4 FILLER_123_239 ();
 FILLCELL_X1 FILLER_123_243 ();
 FILLCELL_X8 FILLER_123_251 ();
 FILLCELL_X4 FILLER_123_263 ();
 FILLCELL_X4 FILLER_123_274 ();
 FILLCELL_X8 FILLER_123_312 ();
 FILLCELL_X1 FILLER_123_320 ();
 FILLCELL_X4 FILLER_123_328 ();
 FILLCELL_X2 FILLER_123_332 ();
 FILLCELL_X1 FILLER_123_334 ();
 FILLCELL_X1 FILLER_123_342 ();
 FILLCELL_X8 FILLER_123_350 ();
 FILLCELL_X4 FILLER_123_365 ();
 FILLCELL_X4 FILLER_123_396 ();
 FILLCELL_X1 FILLER_123_400 ();
 FILLCELL_X1 FILLER_123_405 ();
 FILLCELL_X8 FILLER_123_409 ();
 FILLCELL_X1 FILLER_123_417 ();
 FILLCELL_X8 FILLER_123_459 ();
 FILLCELL_X4 FILLER_123_467 ();
 FILLCELL_X2 FILLER_123_471 ();
 FILLCELL_X1 FILLER_123_473 ();
 FILLCELL_X4 FILLER_123_481 ();
 FILLCELL_X1 FILLER_123_485 ();
 FILLCELL_X16 FILLER_123_513 ();
 FILLCELL_X2 FILLER_123_529 ();
 FILLCELL_X1 FILLER_123_531 ();
 FILLCELL_X16 FILLER_123_539 ();
 FILLCELL_X4 FILLER_123_555 ();
 FILLCELL_X1 FILLER_123_559 ();
 FILLCELL_X1 FILLER_123_594 ();
 FILLCELL_X4 FILLER_123_602 ();
 FILLCELL_X1 FILLER_123_630 ();
 FILLCELL_X16 FILLER_123_652 ();
 FILLCELL_X4 FILLER_123_668 ();
 FILLCELL_X4 FILLER_123_692 ();
 FILLCELL_X1 FILLER_123_696 ();
 FILLCELL_X1 FILLER_123_737 ();
 FILLCELL_X4 FILLER_123_756 ();
 FILLCELL_X8 FILLER_123_780 ();
 FILLCELL_X4 FILLER_123_788 ();
 FILLCELL_X2 FILLER_123_806 ();
 FILLCELL_X1 FILLER_123_808 ();
 FILLCELL_X4 FILLER_123_816 ();
 FILLCELL_X2 FILLER_123_820 ();
 FILLCELL_X2 FILLER_123_854 ();
 FILLCELL_X2 FILLER_123_859 ();
 FILLCELL_X1 FILLER_123_861 ();
 FILLCELL_X1 FILLER_123_869 ();
 FILLCELL_X1 FILLER_123_890 ();
 FILLCELL_X8 FILLER_123_899 ();
 FILLCELL_X4 FILLER_123_907 ();
 FILLCELL_X1 FILLER_123_911 ();
 FILLCELL_X1 FILLER_123_929 ();
 FILLCELL_X1 FILLER_123_954 ();
 FILLCELL_X1 FILLER_123_961 ();
 FILLCELL_X1 FILLER_123_965 ();
 FILLCELL_X2 FILLER_123_977 ();
 FILLCELL_X1 FILLER_123_985 ();
 FILLCELL_X2 FILLER_123_990 ();
 FILLCELL_X1 FILLER_123_996 ();
 FILLCELL_X2 FILLER_123_1019 ();
 FILLCELL_X2 FILLER_123_1057 ();
 FILLCELL_X8 FILLER_123_1062 ();
 FILLCELL_X2 FILLER_123_1083 ();
 FILLCELL_X8 FILLER_123_1088 ();
 FILLCELL_X4 FILLER_123_1096 ();
 FILLCELL_X2 FILLER_123_1100 ();
 FILLCELL_X2 FILLER_123_1140 ();
 FILLCELL_X1 FILLER_123_1149 ();
 FILLCELL_X2 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1177 ();
 FILLCELL_X8 FILLER_123_1209 ();
 FILLCELL_X16 FILLER_123_1220 ();
 FILLCELL_X4 FILLER_123_1236 ();
 FILLCELL_X8 FILLER_123_1243 ();
 FILLCELL_X4 FILLER_123_1251 ();
 FILLCELL_X2 FILLER_124_1 ();
 FILLCELL_X1 FILLER_124_3 ();
 FILLCELL_X4 FILLER_124_24 ();
 FILLCELL_X1 FILLER_124_28 ();
 FILLCELL_X2 FILLER_124_36 ();
 FILLCELL_X2 FILLER_124_48 ();
 FILLCELL_X1 FILLER_124_50 ();
 FILLCELL_X2 FILLER_124_58 ();
 FILLCELL_X1 FILLER_124_60 ();
 FILLCELL_X16 FILLER_124_81 ();
 FILLCELL_X2 FILLER_124_97 ();
 FILLCELL_X8 FILLER_124_123 ();
 FILLCELL_X1 FILLER_124_131 ();
 FILLCELL_X4 FILLER_124_136 ();
 FILLCELL_X16 FILLER_124_155 ();
 FILLCELL_X8 FILLER_124_171 ();
 FILLCELL_X1 FILLER_124_181 ();
 FILLCELL_X2 FILLER_124_207 ();
 FILLCELL_X16 FILLER_124_232 ();
 FILLCELL_X1 FILLER_124_248 ();
 FILLCELL_X2 FILLER_124_256 ();
 FILLCELL_X1 FILLER_124_258 ();
 FILLCELL_X2 FILLER_124_279 ();
 FILLCELL_X4 FILLER_124_308 ();
 FILLCELL_X1 FILLER_124_312 ();
 FILLCELL_X4 FILLER_124_320 ();
 FILLCELL_X1 FILLER_124_371 ();
 FILLCELL_X4 FILLER_124_379 ();
 FILLCELL_X2 FILLER_124_383 ();
 FILLCELL_X1 FILLER_124_385 ();
 FILLCELL_X1 FILLER_124_401 ();
 FILLCELL_X1 FILLER_124_410 ();
 FILLCELL_X2 FILLER_124_414 ();
 FILLCELL_X8 FILLER_124_461 ();
 FILLCELL_X2 FILLER_124_469 ();
 FILLCELL_X1 FILLER_124_471 ();
 FILLCELL_X4 FILLER_124_492 ();
 FILLCELL_X4 FILLER_124_541 ();
 FILLCELL_X2 FILLER_124_545 ();
 FILLCELL_X1 FILLER_124_547 ();
 FILLCELL_X4 FILLER_124_555 ();
 FILLCELL_X2 FILLER_124_559 ();
 FILLCELL_X1 FILLER_124_561 ();
 FILLCELL_X4 FILLER_124_589 ();
 FILLCELL_X2 FILLER_124_593 ();
 FILLCELL_X1 FILLER_124_595 ();
 FILLCELL_X16 FILLER_124_603 ();
 FILLCELL_X1 FILLER_124_619 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X1 FILLER_124_638 ();
 FILLCELL_X2 FILLER_124_648 ();
 FILLCELL_X1 FILLER_124_670 ();
 FILLCELL_X2 FILLER_124_678 ();
 FILLCELL_X16 FILLER_124_687 ();
 FILLCELL_X1 FILLER_124_703 ();
 FILLCELL_X4 FILLER_124_711 ();
 FILLCELL_X1 FILLER_124_715 ();
 FILLCELL_X16 FILLER_124_723 ();
 FILLCELL_X2 FILLER_124_755 ();
 FILLCELL_X8 FILLER_124_771 ();
 FILLCELL_X4 FILLER_124_779 ();
 FILLCELL_X1 FILLER_124_783 ();
 FILLCELL_X16 FILLER_124_818 ();
 FILLCELL_X8 FILLER_124_834 ();
 FILLCELL_X2 FILLER_124_842 ();
 FILLCELL_X4 FILLER_124_848 ();
 FILLCELL_X2 FILLER_124_852 ();
 FILLCELL_X4 FILLER_124_866 ();
 FILLCELL_X2 FILLER_124_877 ();
 FILLCELL_X8 FILLER_124_885 ();
 FILLCELL_X4 FILLER_124_898 ();
 FILLCELL_X1 FILLER_124_902 ();
 FILLCELL_X8 FILLER_124_921 ();
 FILLCELL_X4 FILLER_124_929 ();
 FILLCELL_X1 FILLER_124_933 ();
 FILLCELL_X16 FILLER_124_941 ();
 FILLCELL_X2 FILLER_124_968 ();
 FILLCELL_X4 FILLER_124_973 ();
 FILLCELL_X1 FILLER_124_988 ();
 FILLCELL_X1 FILLER_124_992 ();
 FILLCELL_X8 FILLER_124_1011 ();
 FILLCELL_X4 FILLER_124_1026 ();
 FILLCELL_X8 FILLER_124_1033 ();
 FILLCELL_X2 FILLER_124_1041 ();
 FILLCELL_X4 FILLER_124_1098 ();
 FILLCELL_X2 FILLER_124_1102 ();
 FILLCELL_X2 FILLER_124_1108 ();
 FILLCELL_X2 FILLER_124_1128 ();
 FILLCELL_X1 FILLER_124_1130 ();
 FILLCELL_X1 FILLER_124_1135 ();
 FILLCELL_X1 FILLER_124_1141 ();
 FILLCELL_X1 FILLER_124_1162 ();
 FILLCELL_X16 FILLER_124_1168 ();
 FILLCELL_X32 FILLER_124_1192 ();
 FILLCELL_X16 FILLER_124_1224 ();
 FILLCELL_X8 FILLER_124_1240 ();
 FILLCELL_X4 FILLER_124_1248 ();
 FILLCELL_X2 FILLER_124_1252 ();
 FILLCELL_X1 FILLER_124_1254 ();
 FILLCELL_X16 FILLER_125_1 ();
 FILLCELL_X8 FILLER_125_17 ();
 FILLCELL_X4 FILLER_125_25 ();
 FILLCELL_X2 FILLER_125_29 ();
 FILLCELL_X1 FILLER_125_31 ();
 FILLCELL_X4 FILLER_125_59 ();
 FILLCELL_X1 FILLER_125_63 ();
 FILLCELL_X4 FILLER_125_71 ();
 FILLCELL_X1 FILLER_125_75 ();
 FILLCELL_X2 FILLER_125_90 ();
 FILLCELL_X1 FILLER_125_92 ();
 FILLCELL_X2 FILLER_125_120 ();
 FILLCELL_X1 FILLER_125_122 ();
 FILLCELL_X2 FILLER_125_127 ();
 FILLCELL_X4 FILLER_125_173 ();
 FILLCELL_X2 FILLER_125_177 ();
 FILLCELL_X1 FILLER_125_179 ();
 FILLCELL_X2 FILLER_125_187 ();
 FILLCELL_X1 FILLER_125_189 ();
 FILLCELL_X2 FILLER_125_194 ();
 FILLCELL_X2 FILLER_125_244 ();
 FILLCELL_X1 FILLER_125_246 ();
 FILLCELL_X16 FILLER_125_274 ();
 FILLCELL_X2 FILLER_125_290 ();
 FILLCELL_X1 FILLER_125_292 ();
 FILLCELL_X16 FILLER_125_307 ();
 FILLCELL_X4 FILLER_125_330 ();
 FILLCELL_X1 FILLER_125_334 ();
 FILLCELL_X8 FILLER_125_349 ();
 FILLCELL_X2 FILLER_125_357 ();
 FILLCELL_X2 FILLER_125_373 ();
 FILLCELL_X1 FILLER_125_402 ();
 FILLCELL_X16 FILLER_125_410 ();
 FILLCELL_X2 FILLER_125_426 ();
 FILLCELL_X1 FILLER_125_428 ();
 FILLCELL_X4 FILLER_125_436 ();
 FILLCELL_X1 FILLER_125_440 ();
 FILLCELL_X16 FILLER_125_465 ();
 FILLCELL_X8 FILLER_125_481 ();
 FILLCELL_X1 FILLER_125_489 ();
 FILLCELL_X16 FILLER_125_515 ();
 FILLCELL_X2 FILLER_125_531 ();
 FILLCELL_X2 FILLER_125_560 ();
 FILLCELL_X8 FILLER_125_575 ();
 FILLCELL_X1 FILLER_125_583 ();
 FILLCELL_X4 FILLER_125_604 ();
 FILLCELL_X2 FILLER_125_608 ();
 FILLCELL_X1 FILLER_125_610 ();
 FILLCELL_X2 FILLER_125_631 ();
 FILLCELL_X1 FILLER_125_633 ();
 FILLCELL_X8 FILLER_125_650 ();
 FILLCELL_X2 FILLER_125_658 ();
 FILLCELL_X1 FILLER_125_660 ();
 FILLCELL_X4 FILLER_125_713 ();
 FILLCELL_X2 FILLER_125_717 ();
 FILLCELL_X2 FILLER_125_746 ();
 FILLCELL_X4 FILLER_125_788 ();
 FILLCELL_X8 FILLER_125_799 ();
 FILLCELL_X4 FILLER_125_807 ();
 FILLCELL_X2 FILLER_125_852 ();
 FILLCELL_X2 FILLER_125_872 ();
 FILLCELL_X8 FILLER_125_896 ();
 FILLCELL_X1 FILLER_125_904 ();
 FILLCELL_X1 FILLER_125_957 ();
 FILLCELL_X1 FILLER_125_962 ();
 FILLCELL_X2 FILLER_125_967 ();
 FILLCELL_X1 FILLER_125_969 ();
 FILLCELL_X2 FILLER_125_973 ();
 FILLCELL_X4 FILLER_125_982 ();
 FILLCELL_X1 FILLER_125_986 ();
 FILLCELL_X1 FILLER_125_1035 ();
 FILLCELL_X8 FILLER_125_1043 ();
 FILLCELL_X8 FILLER_125_1055 ();
 FILLCELL_X4 FILLER_125_1063 ();
 FILLCELL_X1 FILLER_125_1067 ();
 FILLCELL_X16 FILLER_125_1071 ();
 FILLCELL_X4 FILLER_125_1097 ();
 FILLCELL_X16 FILLER_125_1128 ();
 FILLCELL_X2 FILLER_125_1144 ();
 FILLCELL_X1 FILLER_125_1146 ();
 FILLCELL_X8 FILLER_125_1154 ();
 FILLCELL_X1 FILLER_125_1162 ();
 FILLCELL_X1 FILLER_125_1165 ();
 FILLCELL_X32 FILLER_125_1170 ();
 FILLCELL_X32 FILLER_125_1202 ();
 FILLCELL_X16 FILLER_125_1234 ();
 FILLCELL_X4 FILLER_125_1250 ();
 FILLCELL_X1 FILLER_125_1254 ();
 FILLCELL_X8 FILLER_126_1 ();
 FILLCELL_X4 FILLER_126_9 ();
 FILLCELL_X1 FILLER_126_13 ();
 FILLCELL_X1 FILLER_126_46 ();
 FILLCELL_X2 FILLER_126_74 ();
 FILLCELL_X8 FILLER_126_90 ();
 FILLCELL_X2 FILLER_126_98 ();
 FILLCELL_X1 FILLER_126_100 ();
 FILLCELL_X2 FILLER_126_108 ();
 FILLCELL_X8 FILLER_126_148 ();
 FILLCELL_X8 FILLER_126_163 ();
 FILLCELL_X4 FILLER_126_171 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X2 FILLER_126_225 ();
 FILLCELL_X1 FILLER_126_227 ();
 FILLCELL_X16 FILLER_126_238 ();
 FILLCELL_X4 FILLER_126_254 ();
 FILLCELL_X2 FILLER_126_258 ();
 FILLCELL_X1 FILLER_126_260 ();
 FILLCELL_X2 FILLER_126_268 ();
 FILLCELL_X8 FILLER_126_311 ();
 FILLCELL_X4 FILLER_126_319 ();
 FILLCELL_X1 FILLER_126_350 ();
 FILLCELL_X16 FILLER_126_372 ();
 FILLCELL_X1 FILLER_126_388 ();
 FILLCELL_X8 FILLER_126_409 ();
 FILLCELL_X4 FILLER_126_417 ();
 FILLCELL_X1 FILLER_126_421 ();
 FILLCELL_X1 FILLER_126_442 ();
 FILLCELL_X2 FILLER_126_481 ();
 FILLCELL_X1 FILLER_126_483 ();
 FILLCELL_X4 FILLER_126_491 ();
 FILLCELL_X1 FILLER_126_502 ();
 FILLCELL_X1 FILLER_126_510 ();
 FILLCELL_X1 FILLER_126_531 ();
 FILLCELL_X1 FILLER_126_539 ();
 FILLCELL_X2 FILLER_126_547 ();
 FILLCELL_X4 FILLER_126_556 ();
 FILLCELL_X1 FILLER_126_560 ();
 FILLCELL_X8 FILLER_126_581 ();
 FILLCELL_X4 FILLER_126_589 ();
 FILLCELL_X2 FILLER_126_593 ();
 FILLCELL_X1 FILLER_126_595 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X4 FILLER_126_632 ();
 FILLCELL_X2 FILLER_126_636 ();
 FILLCELL_X8 FILLER_126_659 ();
 FILLCELL_X4 FILLER_126_667 ();
 FILLCELL_X1 FILLER_126_671 ();
 FILLCELL_X8 FILLER_126_679 ();
 FILLCELL_X2 FILLER_126_687 ();
 FILLCELL_X1 FILLER_126_716 ();
 FILLCELL_X8 FILLER_126_724 ();
 FILLCELL_X4 FILLER_126_732 ();
 FILLCELL_X8 FILLER_126_753 ();
 FILLCELL_X2 FILLER_126_761 ();
 FILLCELL_X1 FILLER_126_809 ();
 FILLCELL_X4 FILLER_126_859 ();
 FILLCELL_X1 FILLER_126_874 ();
 FILLCELL_X2 FILLER_126_909 ();
 FILLCELL_X1 FILLER_126_911 ();
 FILLCELL_X4 FILLER_126_918 ();
 FILLCELL_X2 FILLER_126_942 ();
 FILLCELL_X1 FILLER_126_944 ();
 FILLCELL_X1 FILLER_126_965 ();
 FILLCELL_X4 FILLER_126_981 ();
 FILLCELL_X2 FILLER_126_995 ();
 FILLCELL_X4 FILLER_126_1008 ();
 FILLCELL_X4 FILLER_126_1017 ();
 FILLCELL_X2 FILLER_126_1025 ();
 FILLCELL_X1 FILLER_126_1027 ();
 FILLCELL_X4 FILLER_126_1035 ();
 FILLCELL_X4 FILLER_126_1085 ();
 FILLCELL_X2 FILLER_126_1089 ();
 FILLCELL_X2 FILLER_126_1097 ();
 FILLCELL_X1 FILLER_126_1099 ();
 FILLCELL_X4 FILLER_126_1107 ();
 FILLCELL_X1 FILLER_126_1111 ();
 FILLCELL_X4 FILLER_126_1123 ();
 FILLCELL_X1 FILLER_126_1127 ();
 FILLCELL_X4 FILLER_126_1156 ();
 FILLCELL_X4 FILLER_126_1165 ();
 FILLCELL_X2 FILLER_126_1169 ();
 FILLCELL_X32 FILLER_126_1178 ();
 FILLCELL_X8 FILLER_126_1210 ();
 FILLCELL_X32 FILLER_126_1221 ();
 FILLCELL_X2 FILLER_126_1253 ();
 FILLCELL_X4 FILLER_127_28 ();
 FILLCELL_X2 FILLER_127_32 ();
 FILLCELL_X8 FILLER_127_48 ();
 FILLCELL_X4 FILLER_127_56 ();
 FILLCELL_X2 FILLER_127_60 ();
 FILLCELL_X1 FILLER_127_62 ();
 FILLCELL_X8 FILLER_127_70 ();
 FILLCELL_X4 FILLER_127_78 ();
 FILLCELL_X1 FILLER_127_129 ();
 FILLCELL_X2 FILLER_127_158 ();
 FILLCELL_X4 FILLER_127_180 ();
 FILLCELL_X2 FILLER_127_188 ();
 FILLCELL_X1 FILLER_127_190 ();
 FILLCELL_X8 FILLER_127_195 ();
 FILLCELL_X1 FILLER_127_203 ();
 FILLCELL_X4 FILLER_127_224 ();
 FILLCELL_X1 FILLER_127_228 ();
 FILLCELL_X1 FILLER_127_236 ();
 FILLCELL_X2 FILLER_127_257 ();
 FILLCELL_X1 FILLER_127_259 ();
 FILLCELL_X4 FILLER_127_281 ();
 FILLCELL_X1 FILLER_127_285 ();
 FILLCELL_X4 FILLER_127_300 ();
 FILLCELL_X16 FILLER_127_311 ();
 FILLCELL_X2 FILLER_127_327 ();
 FILLCELL_X2 FILLER_127_336 ();
 FILLCELL_X4 FILLER_127_365 ();
 FILLCELL_X2 FILLER_127_376 ();
 FILLCELL_X8 FILLER_127_380 ();
 FILLCELL_X4 FILLER_127_388 ();
 FILLCELL_X2 FILLER_127_392 ();
 FILLCELL_X8 FILLER_127_401 ();
 FILLCELL_X4 FILLER_127_409 ();
 FILLCELL_X2 FILLER_127_413 ();
 FILLCELL_X1 FILLER_127_415 ();
 FILLCELL_X2 FILLER_127_429 ();
 FILLCELL_X1 FILLER_127_459 ();
 FILLCELL_X2 FILLER_127_474 ();
 FILLCELL_X16 FILLER_127_496 ();
 FILLCELL_X2 FILLER_127_512 ();
 FILLCELL_X2 FILLER_127_518 ();
 FILLCELL_X1 FILLER_127_520 ();
 FILLCELL_X2 FILLER_127_535 ();
 FILLCELL_X8 FILLER_127_544 ();
 FILLCELL_X1 FILLER_127_559 ();
 FILLCELL_X8 FILLER_127_567 ();
 FILLCELL_X4 FILLER_127_575 ();
 FILLCELL_X1 FILLER_127_579 ();
 FILLCELL_X8 FILLER_127_587 ();
 FILLCELL_X4 FILLER_127_595 ();
 FILLCELL_X2 FILLER_127_599 ();
 FILLCELL_X16 FILLER_127_615 ();
 FILLCELL_X2 FILLER_127_631 ();
 FILLCELL_X8 FILLER_127_660 ();
 FILLCELL_X2 FILLER_127_668 ();
 FILLCELL_X2 FILLER_127_678 ();
 FILLCELL_X4 FILLER_127_692 ();
 FILLCELL_X1 FILLER_127_696 ();
 FILLCELL_X2 FILLER_127_702 ();
 FILLCELL_X1 FILLER_127_704 ();
 FILLCELL_X1 FILLER_127_712 ();
 FILLCELL_X2 FILLER_127_720 ();
 FILLCELL_X4 FILLER_127_732 ();
 FILLCELL_X2 FILLER_127_736 ();
 FILLCELL_X1 FILLER_127_738 ();
 FILLCELL_X4 FILLER_127_753 ();
 FILLCELL_X2 FILLER_127_757 ();
 FILLCELL_X1 FILLER_127_759 ();
 FILLCELL_X16 FILLER_127_774 ();
 FILLCELL_X1 FILLER_127_831 ();
 FILLCELL_X2 FILLER_127_849 ();
 FILLCELL_X1 FILLER_127_851 ();
 FILLCELL_X4 FILLER_127_862 ();
 FILLCELL_X1 FILLER_127_884 ();
 FILLCELL_X2 FILLER_127_899 ();
 FILLCELL_X2 FILLER_127_918 ();
 FILLCELL_X1 FILLER_127_929 ();
 FILLCELL_X1 FILLER_127_941 ();
 FILLCELL_X2 FILLER_127_968 ();
 FILLCELL_X1 FILLER_127_970 ();
 FILLCELL_X1 FILLER_127_978 ();
 FILLCELL_X1 FILLER_127_990 ();
 FILLCELL_X1 FILLER_127_995 ();
 FILLCELL_X2 FILLER_127_999 ();
 FILLCELL_X2 FILLER_127_1008 ();
 FILLCELL_X8 FILLER_127_1013 ();
 FILLCELL_X1 FILLER_127_1021 ();
 FILLCELL_X8 FILLER_127_1047 ();
 FILLCELL_X4 FILLER_127_1055 ();
 FILLCELL_X1 FILLER_127_1059 ();
 FILLCELL_X4 FILLER_127_1069 ();
 FILLCELL_X2 FILLER_127_1073 ();
 FILLCELL_X2 FILLER_127_1103 ();
 FILLCELL_X1 FILLER_127_1170 ();
 FILLCELL_X32 FILLER_127_1191 ();
 FILLCELL_X16 FILLER_127_1223 ();
 FILLCELL_X8 FILLER_127_1239 ();
 FILLCELL_X2 FILLER_127_1247 ();
 FILLCELL_X1 FILLER_127_1249 ();
 FILLCELL_X2 FILLER_127_1253 ();
 FILLCELL_X4 FILLER_128_28 ();
 FILLCELL_X2 FILLER_128_32 ();
 FILLCELL_X1 FILLER_128_34 ();
 FILLCELL_X8 FILLER_128_56 ();
 FILLCELL_X4 FILLER_128_64 ();
 FILLCELL_X2 FILLER_128_68 ();
 FILLCELL_X1 FILLER_128_70 ();
 FILLCELL_X2 FILLER_128_78 ();
 FILLCELL_X1 FILLER_128_80 ();
 FILLCELL_X4 FILLER_128_88 ();
 FILLCELL_X2 FILLER_128_92 ();
 FILLCELL_X4 FILLER_128_101 ();
 FILLCELL_X2 FILLER_128_105 ();
 FILLCELL_X4 FILLER_128_127 ();
 FILLCELL_X4 FILLER_128_145 ();
 FILLCELL_X1 FILLER_128_149 ();
 FILLCELL_X4 FILLER_128_167 ();
 FILLCELL_X4 FILLER_128_205 ();
 FILLCELL_X1 FILLER_128_209 ();
 FILLCELL_X2 FILLER_128_217 ();
 FILLCELL_X4 FILLER_128_233 ();
 FILLCELL_X1 FILLER_128_237 ();
 FILLCELL_X4 FILLER_128_247 ();
 FILLCELL_X1 FILLER_128_251 ();
 FILLCELL_X1 FILLER_128_262 ();
 FILLCELL_X2 FILLER_128_277 ();
 FILLCELL_X8 FILLER_128_316 ();
 FILLCELL_X2 FILLER_128_324 ();
 FILLCELL_X4 FILLER_128_351 ();
 FILLCELL_X2 FILLER_128_355 ();
 FILLCELL_X1 FILLER_128_357 ();
 FILLCELL_X2 FILLER_128_365 ();
 FILLCELL_X4 FILLER_128_415 ();
 FILLCELL_X1 FILLER_128_444 ();
 FILLCELL_X8 FILLER_128_452 ();
 FILLCELL_X2 FILLER_128_460 ();
 FILLCELL_X1 FILLER_128_462 ();
 FILLCELL_X1 FILLER_128_468 ();
 FILLCELL_X4 FILLER_128_476 ();
 FILLCELL_X1 FILLER_128_480 ();
 FILLCELL_X2 FILLER_128_488 ();
 FILLCELL_X2 FILLER_128_517 ();
 FILLCELL_X1 FILLER_128_519 ();
 FILLCELL_X1 FILLER_128_547 ();
 FILLCELL_X4 FILLER_128_555 ();
 FILLCELL_X1 FILLER_128_566 ();
 FILLCELL_X4 FILLER_128_574 ();
 FILLCELL_X2 FILLER_128_578 ();
 FILLCELL_X8 FILLER_128_583 ();
 FILLCELL_X4 FILLER_128_591 ();
 FILLCELL_X1 FILLER_128_595 ();
 FILLCELL_X2 FILLER_128_612 ();
 FILLCELL_X1 FILLER_128_614 ();
 FILLCELL_X2 FILLER_128_632 ();
 FILLCELL_X1 FILLER_128_634 ();
 FILLCELL_X4 FILLER_128_642 ();
 FILLCELL_X1 FILLER_128_646 ();
 FILLCELL_X2 FILLER_128_687 ();
 FILLCELL_X1 FILLER_128_689 ();
 FILLCELL_X16 FILLER_128_697 ();
 FILLCELL_X4 FILLER_128_727 ();
 FILLCELL_X1 FILLER_128_731 ();
 FILLCELL_X2 FILLER_128_746 ();
 FILLCELL_X16 FILLER_128_775 ();
 FILLCELL_X8 FILLER_128_791 ();
 FILLCELL_X2 FILLER_128_799 ();
 FILLCELL_X2 FILLER_128_815 ();
 FILLCELL_X2 FILLER_128_831 ();
 FILLCELL_X2 FILLER_128_852 ();
 FILLCELL_X1 FILLER_128_854 ();
 FILLCELL_X2 FILLER_128_874 ();
 FILLCELL_X1 FILLER_128_876 ();
 FILLCELL_X2 FILLER_128_901 ();
 FILLCELL_X1 FILLER_128_903 ();
 FILLCELL_X2 FILLER_128_915 ();
 FILLCELL_X2 FILLER_128_926 ();
 FILLCELL_X4 FILLER_128_965 ();
 FILLCELL_X2 FILLER_128_969 ();
 FILLCELL_X1 FILLER_128_971 ();
 FILLCELL_X4 FILLER_128_996 ();
 FILLCELL_X2 FILLER_128_1011 ();
 FILLCELL_X1 FILLER_128_1013 ();
 FILLCELL_X4 FILLER_128_1017 ();
 FILLCELL_X2 FILLER_128_1021 ();
 FILLCELL_X4 FILLER_128_1030 ();
 FILLCELL_X8 FILLER_128_1037 ();
 FILLCELL_X2 FILLER_128_1045 ();
 FILLCELL_X4 FILLER_128_1058 ();
 FILLCELL_X1 FILLER_128_1079 ();
 FILLCELL_X8 FILLER_128_1090 ();
 FILLCELL_X2 FILLER_128_1098 ();
 FILLCELL_X16 FILLER_128_1110 ();
 FILLCELL_X1 FILLER_128_1126 ();
 FILLCELL_X4 FILLER_128_1130 ();
 FILLCELL_X1 FILLER_128_1134 ();
 FILLCELL_X1 FILLER_128_1139 ();
 FILLCELL_X4 FILLER_128_1146 ();
 FILLCELL_X4 FILLER_128_1153 ();
 FILLCELL_X1 FILLER_128_1157 ();
 FILLCELL_X4 FILLER_128_1164 ();
 FILLCELL_X32 FILLER_128_1172 ();
 FILLCELL_X16 FILLER_128_1204 ();
 FILLCELL_X4 FILLER_128_1220 ();
 FILLCELL_X2 FILLER_128_1224 ();
 FILLCELL_X16 FILLER_128_1229 ();
 FILLCELL_X8 FILLER_128_1245 ();
 FILLCELL_X2 FILLER_128_1253 ();
 FILLCELL_X16 FILLER_129_1 ();
 FILLCELL_X4 FILLER_129_51 ();
 FILLCELL_X1 FILLER_129_55 ();
 FILLCELL_X2 FILLER_129_76 ();
 FILLCELL_X16 FILLER_129_99 ();
 FILLCELL_X4 FILLER_129_115 ();
 FILLCELL_X1 FILLER_129_139 ();
 FILLCELL_X16 FILLER_129_161 ();
 FILLCELL_X8 FILLER_129_177 ();
 FILLCELL_X8 FILLER_129_206 ();
 FILLCELL_X1 FILLER_129_234 ();
 FILLCELL_X1 FILLER_129_239 ();
 FILLCELL_X1 FILLER_129_269 ();
 FILLCELL_X2 FILLER_129_295 ();
 FILLCELL_X1 FILLER_129_301 ();
 FILLCELL_X4 FILLER_129_329 ();
 FILLCELL_X2 FILLER_129_333 ();
 FILLCELL_X1 FILLER_129_335 ();
 FILLCELL_X8 FILLER_129_370 ();
 FILLCELL_X4 FILLER_129_378 ();
 FILLCELL_X1 FILLER_129_382 ();
 FILLCELL_X4 FILLER_129_405 ();
 FILLCELL_X1 FILLER_129_409 ();
 FILLCELL_X2 FILLER_129_457 ();
 FILLCELL_X1 FILLER_129_459 ();
 FILLCELL_X4 FILLER_129_485 ();
 FILLCELL_X2 FILLER_129_520 ();
 FILLCELL_X1 FILLER_129_522 ();
 FILLCELL_X4 FILLER_129_530 ();
 FILLCELL_X1 FILLER_129_534 ();
 FILLCELL_X4 FILLER_129_542 ();
 FILLCELL_X1 FILLER_129_546 ();
 FILLCELL_X4 FILLER_129_567 ();
 FILLCELL_X4 FILLER_129_594 ();
 FILLCELL_X2 FILLER_129_598 ();
 FILLCELL_X1 FILLER_129_600 ();
 FILLCELL_X2 FILLER_129_615 ();
 FILLCELL_X1 FILLER_129_617 ();
 FILLCELL_X4 FILLER_129_632 ();
 FILLCELL_X16 FILLER_129_647 ();
 FILLCELL_X4 FILLER_129_670 ();
 FILLCELL_X2 FILLER_129_674 ();
 FILLCELL_X4 FILLER_129_683 ();
 FILLCELL_X1 FILLER_129_687 ();
 FILLCELL_X16 FILLER_129_695 ();
 FILLCELL_X2 FILLER_129_711 ();
 FILLCELL_X1 FILLER_129_745 ();
 FILLCELL_X1 FILLER_129_751 ();
 FILLCELL_X1 FILLER_129_792 ();
 FILLCELL_X1 FILLER_129_830 ();
 FILLCELL_X4 FILLER_129_849 ();
 FILLCELL_X2 FILLER_129_853 ();
 FILLCELL_X1 FILLER_129_877 ();
 FILLCELL_X2 FILLER_129_893 ();
 FILLCELL_X1 FILLER_129_895 ();
 FILLCELL_X4 FILLER_129_909 ();
 FILLCELL_X4 FILLER_129_916 ();
 FILLCELL_X2 FILLER_129_927 ();
 FILLCELL_X4 FILLER_129_941 ();
 FILLCELL_X1 FILLER_129_945 ();
 FILLCELL_X2 FILLER_129_949 ();
 FILLCELL_X1 FILLER_129_951 ();
 FILLCELL_X2 FILLER_129_955 ();
 FILLCELL_X1 FILLER_129_957 ();
 FILLCELL_X8 FILLER_129_971 ();
 FILLCELL_X2 FILLER_129_994 ();
 FILLCELL_X1 FILLER_129_1014 ();
 FILLCELL_X2 FILLER_129_1024 ();
 FILLCELL_X2 FILLER_129_1029 ();
 FILLCELL_X1 FILLER_129_1031 ();
 FILLCELL_X4 FILLER_129_1052 ();
 FILLCELL_X8 FILLER_129_1068 ();
 FILLCELL_X2 FILLER_129_1076 ();
 FILLCELL_X2 FILLER_129_1083 ();
 FILLCELL_X1 FILLER_129_1085 ();
 FILLCELL_X4 FILLER_129_1118 ();
 FILLCELL_X2 FILLER_129_1122 ();
 FILLCELL_X4 FILLER_129_1144 ();
 FILLCELL_X2 FILLER_129_1148 ();
 FILLCELL_X2 FILLER_129_1152 ();
 FILLCELL_X4 FILLER_129_1163 ();
 FILLCELL_X32 FILLER_129_1174 ();
 FILLCELL_X8 FILLER_129_1206 ();
 FILLCELL_X2 FILLER_129_1214 ();
 FILLCELL_X1 FILLER_129_1216 ();
 FILLCELL_X16 FILLER_129_1220 ();
 FILLCELL_X8 FILLER_129_1236 ();
 FILLCELL_X4 FILLER_129_1244 ();
 FILLCELL_X1 FILLER_129_1248 ();
 FILLCELL_X2 FILLER_129_1252 ();
 FILLCELL_X1 FILLER_129_1254 ();
 FILLCELL_X8 FILLER_130_1 ();
 FILLCELL_X2 FILLER_130_9 ();
 FILLCELL_X4 FILLER_130_19 ();
 FILLCELL_X2 FILLER_130_23 ();
 FILLCELL_X1 FILLER_130_25 ();
 FILLCELL_X4 FILLER_130_40 ();
 FILLCELL_X1 FILLER_130_44 ();
 FILLCELL_X2 FILLER_130_52 ();
 FILLCELL_X1 FILLER_130_54 ();
 FILLCELL_X4 FILLER_130_75 ();
 FILLCELL_X1 FILLER_130_79 ();
 FILLCELL_X4 FILLER_130_87 ();
 FILLCELL_X1 FILLER_130_91 ();
 FILLCELL_X4 FILLER_130_112 ();
 FILLCELL_X16 FILLER_130_123 ();
 FILLCELL_X8 FILLER_130_139 ();
 FILLCELL_X2 FILLER_130_147 ();
 FILLCELL_X8 FILLER_130_156 ();
 FILLCELL_X4 FILLER_130_164 ();
 FILLCELL_X1 FILLER_130_188 ();
 FILLCELL_X2 FILLER_130_196 ();
 FILLCELL_X1 FILLER_130_205 ();
 FILLCELL_X2 FILLER_130_213 ();
 FILLCELL_X2 FILLER_130_222 ();
 FILLCELL_X1 FILLER_130_224 ();
 FILLCELL_X4 FILLER_130_232 ();
 FILLCELL_X2 FILLER_130_236 ();
 FILLCELL_X1 FILLER_130_238 ();
 FILLCELL_X2 FILLER_130_256 ();
 FILLCELL_X1 FILLER_130_258 ();
 FILLCELL_X8 FILLER_130_266 ();
 FILLCELL_X2 FILLER_130_274 ();
 FILLCELL_X4 FILLER_130_303 ();
 FILLCELL_X1 FILLER_130_307 ();
 FILLCELL_X1 FILLER_130_315 ();
 FILLCELL_X2 FILLER_130_323 ();
 FILLCELL_X1 FILLER_130_392 ();
 FILLCELL_X8 FILLER_130_395 ();
 FILLCELL_X2 FILLER_130_403 ();
 FILLCELL_X1 FILLER_130_405 ();
 FILLCELL_X4 FILLER_130_448 ();
 FILLCELL_X2 FILLER_130_452 ();
 FILLCELL_X1 FILLER_130_481 ();
 FILLCELL_X8 FILLER_130_496 ();
 FILLCELL_X1 FILLER_130_504 ();
 FILLCELL_X16 FILLER_130_532 ();
 FILLCELL_X8 FILLER_130_548 ();
 FILLCELL_X4 FILLER_130_556 ();
 FILLCELL_X1 FILLER_130_560 ();
 FILLCELL_X8 FILLER_130_591 ();
 FILLCELL_X2 FILLER_130_599 ();
 FILLCELL_X2 FILLER_130_614 ();
 FILLCELL_X1 FILLER_130_616 ();
 FILLCELL_X1 FILLER_130_632 ();
 FILLCELL_X4 FILLER_130_663 ();
 FILLCELL_X2 FILLER_130_667 ();
 FILLCELL_X1 FILLER_130_669 ();
 FILLCELL_X4 FILLER_130_724 ();
 FILLCELL_X1 FILLER_130_748 ();
 FILLCELL_X2 FILLER_130_763 ();
 FILLCELL_X1 FILLER_130_765 ();
 FILLCELL_X1 FILLER_130_770 ();
 FILLCELL_X1 FILLER_130_783 ();
 FILLCELL_X8 FILLER_130_798 ();
 FILLCELL_X1 FILLER_130_806 ();
 FILLCELL_X8 FILLER_130_821 ();
 FILLCELL_X1 FILLER_130_829 ();
 FILLCELL_X1 FILLER_130_833 ();
 FILLCELL_X2 FILLER_130_860 ();
 FILLCELL_X1 FILLER_130_866 ();
 FILLCELL_X2 FILLER_130_882 ();
 FILLCELL_X1 FILLER_130_884 ();
 FILLCELL_X1 FILLER_130_892 ();
 FILLCELL_X1 FILLER_130_897 ();
 FILLCELL_X1 FILLER_130_905 ();
 FILLCELL_X1 FILLER_130_913 ();
 FILLCELL_X4 FILLER_130_928 ();
 FILLCELL_X2 FILLER_130_932 ();
 FILLCELL_X1 FILLER_130_934 ();
 FILLCELL_X4 FILLER_130_938 ();
 FILLCELL_X4 FILLER_130_944 ();
 FILLCELL_X2 FILLER_130_948 ();
 FILLCELL_X1 FILLER_130_950 ();
 FILLCELL_X4 FILLER_130_957 ();
 FILLCELL_X1 FILLER_130_961 ();
 FILLCELL_X1 FILLER_130_966 ();
 FILLCELL_X8 FILLER_130_974 ();
 FILLCELL_X2 FILLER_130_982 ();
 FILLCELL_X1 FILLER_130_999 ();
 FILLCELL_X1 FILLER_130_1007 ();
 FILLCELL_X2 FILLER_130_1011 ();
 FILLCELL_X1 FILLER_130_1013 ();
 FILLCELL_X1 FILLER_130_1021 ();
 FILLCELL_X8 FILLER_130_1029 ();
 FILLCELL_X8 FILLER_130_1050 ();
 FILLCELL_X2 FILLER_130_1058 ();
 FILLCELL_X2 FILLER_130_1090 ();
 FILLCELL_X1 FILLER_130_1092 ();
 FILLCELL_X2 FILLER_130_1103 ();
 FILLCELL_X8 FILLER_130_1115 ();
 FILLCELL_X2 FILLER_130_1123 ();
 FILLCELL_X1 FILLER_130_1125 ();
 FILLCELL_X2 FILLER_130_1130 ();
 FILLCELL_X1 FILLER_130_1139 ();
 FILLCELL_X32 FILLER_130_1184 ();
 FILLCELL_X8 FILLER_130_1216 ();
 FILLCELL_X4 FILLER_130_1227 ();
 FILLCELL_X1 FILLER_130_1231 ();
 FILLCELL_X16 FILLER_130_1235 ();
 FILLCELL_X4 FILLER_130_1251 ();
 FILLCELL_X4 FILLER_131_28 ();
 FILLCELL_X8 FILLER_131_53 ();
 FILLCELL_X2 FILLER_131_61 ();
 FILLCELL_X4 FILLER_131_70 ();
 FILLCELL_X2 FILLER_131_74 ();
 FILLCELL_X1 FILLER_131_76 ();
 FILLCELL_X2 FILLER_131_84 ();
 FILLCELL_X1 FILLER_131_93 ();
 FILLCELL_X2 FILLER_131_135 ();
 FILLCELL_X1 FILLER_131_164 ();
 FILLCELL_X4 FILLER_131_220 ();
 FILLCELL_X2 FILLER_131_224 ();
 FILLCELL_X2 FILLER_131_246 ();
 FILLCELL_X1 FILLER_131_248 ();
 FILLCELL_X32 FILLER_131_252 ();
 FILLCELL_X4 FILLER_131_284 ();
 FILLCELL_X2 FILLER_131_288 ();
 FILLCELL_X2 FILLER_131_308 ();
 FILLCELL_X8 FILLER_131_326 ();
 FILLCELL_X2 FILLER_131_334 ();
 FILLCELL_X1 FILLER_131_336 ();
 FILLCELL_X16 FILLER_131_344 ();
 FILLCELL_X1 FILLER_131_360 ();
 FILLCELL_X8 FILLER_131_368 ();
 FILLCELL_X4 FILLER_131_383 ();
 FILLCELL_X2 FILLER_131_387 ();
 FILLCELL_X1 FILLER_131_389 ();
 FILLCELL_X8 FILLER_131_393 ();
 FILLCELL_X1 FILLER_131_401 ();
 FILLCELL_X4 FILLER_131_412 ();
 FILLCELL_X1 FILLER_131_416 ();
 FILLCELL_X1 FILLER_131_432 ();
 FILLCELL_X4 FILLER_131_436 ();
 FILLCELL_X2 FILLER_131_481 ();
 FILLCELL_X4 FILLER_131_500 ();
 FILLCELL_X2 FILLER_131_504 ();
 FILLCELL_X1 FILLER_131_506 ();
 FILLCELL_X4 FILLER_131_535 ();
 FILLCELL_X4 FILLER_131_556 ();
 FILLCELL_X2 FILLER_131_560 ();
 FILLCELL_X1 FILLER_131_562 ();
 FILLCELL_X4 FILLER_131_583 ();
 FILLCELL_X2 FILLER_131_587 ();
 FILLCELL_X1 FILLER_131_589 ();
 FILLCELL_X8 FILLER_131_606 ();
 FILLCELL_X2 FILLER_131_630 ();
 FILLCELL_X8 FILLER_131_646 ();
 FILLCELL_X2 FILLER_131_654 ();
 FILLCELL_X4 FILLER_131_683 ();
 FILLCELL_X4 FILLER_131_708 ();
 FILLCELL_X1 FILLER_131_712 ();
 FILLCELL_X2 FILLER_131_720 ();
 FILLCELL_X1 FILLER_131_736 ();
 FILLCELL_X8 FILLER_131_740 ();
 FILLCELL_X4 FILLER_131_748 ();
 FILLCELL_X1 FILLER_131_752 ();
 FILLCELL_X16 FILLER_131_780 ();
 FILLCELL_X1 FILLER_131_810 ();
 FILLCELL_X4 FILLER_131_825 ();
 FILLCELL_X1 FILLER_131_829 ();
 FILLCELL_X2 FILLER_131_845 ();
 FILLCELL_X1 FILLER_131_863 ();
 FILLCELL_X4 FILLER_131_873 ();
 FILLCELL_X2 FILLER_131_909 ();
 FILLCELL_X4 FILLER_131_926 ();
 FILLCELL_X2 FILLER_131_956 ();
 FILLCELL_X1 FILLER_131_958 ();
 FILLCELL_X2 FILLER_131_977 ();
 FILLCELL_X1 FILLER_131_979 ();
 FILLCELL_X2 FILLER_131_985 ();
 FILLCELL_X8 FILLER_131_1000 ();
 FILLCELL_X4 FILLER_131_1015 ();
 FILLCELL_X1 FILLER_131_1019 ();
 FILLCELL_X4 FILLER_131_1025 ();
 FILLCELL_X2 FILLER_131_1029 ();
 FILLCELL_X4 FILLER_131_1049 ();
 FILLCELL_X1 FILLER_131_1053 ();
 FILLCELL_X2 FILLER_131_1059 ();
 FILLCELL_X2 FILLER_131_1076 ();
 FILLCELL_X4 FILLER_131_1154 ();
 FILLCELL_X2 FILLER_131_1158 ();
 FILLCELL_X1 FILLER_131_1165 ();
 FILLCELL_X32 FILLER_131_1179 ();
 FILLCELL_X4 FILLER_131_1211 ();
 FILLCELL_X2 FILLER_131_1215 ();
 FILLCELL_X1 FILLER_131_1217 ();
 FILLCELL_X32 FILLER_131_1221 ();
 FILLCELL_X2 FILLER_131_1253 ();
 FILLCELL_X8 FILLER_132_1 ();
 FILLCELL_X4 FILLER_132_9 ();
 FILLCELL_X4 FILLER_132_40 ();
 FILLCELL_X8 FILLER_132_51 ();
 FILLCELL_X2 FILLER_132_59 ();
 FILLCELL_X8 FILLER_132_88 ();
 FILLCELL_X4 FILLER_132_96 ();
 FILLCELL_X4 FILLER_132_119 ();
 FILLCELL_X2 FILLER_132_123 ();
 FILLCELL_X1 FILLER_132_157 ();
 FILLCELL_X16 FILLER_132_163 ();
 FILLCELL_X2 FILLER_132_179 ();
 FILLCELL_X1 FILLER_132_181 ();
 FILLCELL_X2 FILLER_132_193 ();
 FILLCELL_X1 FILLER_132_195 ();
 FILLCELL_X2 FILLER_132_200 ();
 FILLCELL_X8 FILLER_132_205 ();
 FILLCELL_X4 FILLER_132_213 ();
 FILLCELL_X1 FILLER_132_217 ();
 FILLCELL_X4 FILLER_132_225 ();
 FILLCELL_X1 FILLER_132_229 ();
 FILLCELL_X8 FILLER_132_277 ();
 FILLCELL_X4 FILLER_132_285 ();
 FILLCELL_X2 FILLER_132_289 ();
 FILLCELL_X1 FILLER_132_291 ();
 FILLCELL_X1 FILLER_132_299 ();
 FILLCELL_X2 FILLER_132_310 ();
 FILLCELL_X1 FILLER_132_312 ();
 FILLCELL_X8 FILLER_132_320 ();
 FILLCELL_X2 FILLER_132_328 ();
 FILLCELL_X1 FILLER_132_330 ();
 FILLCELL_X2 FILLER_132_338 ();
 FILLCELL_X1 FILLER_132_340 ();
 FILLCELL_X2 FILLER_132_368 ();
 FILLCELL_X1 FILLER_132_370 ();
 FILLCELL_X4 FILLER_132_378 ();
 FILLCELL_X2 FILLER_132_393 ();
 FILLCELL_X1 FILLER_132_400 ();
 FILLCELL_X4 FILLER_132_410 ();
 FILLCELL_X2 FILLER_132_414 ();
 FILLCELL_X1 FILLER_132_416 ();
 FILLCELL_X2 FILLER_132_424 ();
 FILLCELL_X1 FILLER_132_426 ();
 FILLCELL_X1 FILLER_132_431 ();
 FILLCELL_X2 FILLER_132_444 ();
 FILLCELL_X1 FILLER_132_471 ();
 FILLCELL_X2 FILLER_132_479 ();
 FILLCELL_X2 FILLER_132_495 ();
 FILLCELL_X2 FILLER_132_517 ();
 FILLCELL_X4 FILLER_132_526 ();
 FILLCELL_X1 FILLER_132_530 ();
 FILLCELL_X4 FILLER_132_558 ();
 FILLCELL_X2 FILLER_132_562 ();
 FILLCELL_X1 FILLER_132_564 ();
 FILLCELL_X8 FILLER_132_578 ();
 FILLCELL_X2 FILLER_132_596 ();
 FILLCELL_X4 FILLER_132_616 ();
 FILLCELL_X2 FILLER_132_620 ();
 FILLCELL_X2 FILLER_132_653 ();
 FILLCELL_X1 FILLER_132_655 ();
 FILLCELL_X1 FILLER_132_675 ();
 FILLCELL_X2 FILLER_132_683 ();
 FILLCELL_X2 FILLER_132_692 ();
 FILLCELL_X1 FILLER_132_694 ();
 FILLCELL_X2 FILLER_132_702 ();
 FILLCELL_X1 FILLER_132_704 ();
 FILLCELL_X2 FILLER_132_710 ();
 FILLCELL_X8 FILLER_132_740 ();
 FILLCELL_X2 FILLER_132_748 ();
 FILLCELL_X1 FILLER_132_750 ();
 FILLCELL_X8 FILLER_132_758 ();
 FILLCELL_X1 FILLER_132_766 ();
 FILLCELL_X4 FILLER_132_774 ();
 FILLCELL_X1 FILLER_132_778 ();
 FILLCELL_X1 FILLER_132_799 ();
 FILLCELL_X1 FILLER_132_817 ();
 FILLCELL_X4 FILLER_132_827 ();
 FILLCELL_X2 FILLER_132_831 ();
 FILLCELL_X1 FILLER_132_833 ();
 FILLCELL_X2 FILLER_132_837 ();
 FILLCELL_X1 FILLER_132_846 ();
 FILLCELL_X8 FILLER_132_852 ();
 FILLCELL_X1 FILLER_132_891 ();
 FILLCELL_X1 FILLER_132_894 ();
 FILLCELL_X8 FILLER_132_902 ();
 FILLCELL_X1 FILLER_132_910 ();
 FILLCELL_X1 FILLER_132_920 ();
 FILLCELL_X16 FILLER_132_926 ();
 FILLCELL_X4 FILLER_132_942 ();
 FILLCELL_X1 FILLER_132_946 ();
 FILLCELL_X16 FILLER_132_952 ();
 FILLCELL_X4 FILLER_132_968 ();
 FILLCELL_X1 FILLER_132_972 ();
 FILLCELL_X4 FILLER_132_976 ();
 FILLCELL_X1 FILLER_132_980 ();
 FILLCELL_X4 FILLER_132_1023 ();
 FILLCELL_X1 FILLER_132_1027 ();
 FILLCELL_X2 FILLER_132_1035 ();
 FILLCELL_X16 FILLER_132_1044 ();
 FILLCELL_X1 FILLER_132_1060 ();
 FILLCELL_X1 FILLER_132_1086 ();
 FILLCELL_X1 FILLER_132_1091 ();
 FILLCELL_X4 FILLER_132_1095 ();
 FILLCELL_X2 FILLER_132_1099 ();
 FILLCELL_X1 FILLER_132_1101 ();
 FILLCELL_X4 FILLER_132_1109 ();
 FILLCELL_X2 FILLER_132_1113 ();
 FILLCELL_X1 FILLER_132_1115 ();
 FILLCELL_X4 FILLER_132_1118 ();
 FILLCELL_X1 FILLER_132_1122 ();
 FILLCELL_X2 FILLER_132_1143 ();
 FILLCELL_X2 FILLER_132_1169 ();
 FILLCELL_X32 FILLER_132_1193 ();
 FILLCELL_X1 FILLER_132_1225 ();
 FILLCELL_X8 FILLER_132_1229 ();
 FILLCELL_X8 FILLER_132_1243 ();
 FILLCELL_X4 FILLER_132_1251 ();
 FILLCELL_X16 FILLER_133_1 ();
 FILLCELL_X2 FILLER_133_17 ();
 FILLCELL_X1 FILLER_133_19 ();
 FILLCELL_X2 FILLER_133_92 ();
 FILLCELL_X2 FILLER_133_114 ();
 FILLCELL_X16 FILLER_133_123 ();
 FILLCELL_X2 FILLER_133_139 ();
 FILLCELL_X1 FILLER_133_141 ();
 FILLCELL_X4 FILLER_133_169 ();
 FILLCELL_X2 FILLER_133_173 ();
 FILLCELL_X4 FILLER_133_186 ();
 FILLCELL_X1 FILLER_133_194 ();
 FILLCELL_X8 FILLER_133_257 ();
 FILLCELL_X1 FILLER_133_265 ();
 FILLCELL_X1 FILLER_133_280 ();
 FILLCELL_X4 FILLER_133_301 ();
 FILLCELL_X4 FILLER_133_319 ();
 FILLCELL_X1 FILLER_133_323 ();
 FILLCELL_X16 FILLER_133_337 ();
 FILLCELL_X4 FILLER_133_353 ();
 FILLCELL_X2 FILLER_133_357 ();
 FILLCELL_X2 FILLER_133_386 ();
 FILLCELL_X2 FILLER_133_395 ();
 FILLCELL_X1 FILLER_133_397 ();
 FILLCELL_X1 FILLER_133_402 ();
 FILLCELL_X2 FILLER_133_410 ();
 FILLCELL_X2 FILLER_133_419 ();
 FILLCELL_X2 FILLER_133_428 ();
 FILLCELL_X2 FILLER_133_487 ();
 FILLCELL_X8 FILLER_133_492 ();
 FILLCELL_X2 FILLER_133_500 ();
 FILLCELL_X1 FILLER_133_502 ();
 FILLCELL_X2 FILLER_133_515 ();
 FILLCELL_X32 FILLER_133_544 ();
 FILLCELL_X8 FILLER_133_576 ();
 FILLCELL_X2 FILLER_133_584 ();
 FILLCELL_X1 FILLER_133_586 ();
 FILLCELL_X2 FILLER_133_601 ();
 FILLCELL_X16 FILLER_133_606 ();
 FILLCELL_X4 FILLER_133_622 ();
 FILLCELL_X2 FILLER_133_626 ();
 FILLCELL_X1 FILLER_133_628 ();
 FILLCELL_X4 FILLER_133_652 ();
 FILLCELL_X1 FILLER_133_656 ();
 FILLCELL_X4 FILLER_133_660 ();
 FILLCELL_X2 FILLER_133_664 ();
 FILLCELL_X2 FILLER_133_693 ();
 FILLCELL_X1 FILLER_133_695 ();
 FILLCELL_X8 FILLER_133_728 ();
 FILLCELL_X2 FILLER_133_763 ();
 FILLCELL_X2 FILLER_133_772 ();
 FILLCELL_X1 FILLER_133_774 ();
 FILLCELL_X2 FILLER_133_782 ();
 FILLCELL_X4 FILLER_133_804 ();
 FILLCELL_X2 FILLER_133_808 ();
 FILLCELL_X1 FILLER_133_810 ();
 FILLCELL_X2 FILLER_133_828 ();
 FILLCELL_X4 FILLER_133_842 ();
 FILLCELL_X2 FILLER_133_846 ();
 FILLCELL_X2 FILLER_133_852 ();
 FILLCELL_X16 FILLER_133_863 ();
 FILLCELL_X1 FILLER_133_879 ();
 FILLCELL_X2 FILLER_133_887 ();
 FILLCELL_X1 FILLER_133_889 ();
 FILLCELL_X1 FILLER_133_902 ();
 FILLCELL_X4 FILLER_133_907 ();
 FILLCELL_X1 FILLER_133_911 ();
 FILLCELL_X2 FILLER_133_917 ();
 FILLCELL_X1 FILLER_133_919 ();
 FILLCELL_X1 FILLER_133_944 ();
 FILLCELL_X8 FILLER_133_978 ();
 FILLCELL_X2 FILLER_133_986 ();
 FILLCELL_X1 FILLER_133_988 ();
 FILLCELL_X8 FILLER_133_1005 ();
 FILLCELL_X4 FILLER_133_1013 ();
 FILLCELL_X1 FILLER_133_1017 ();
 FILLCELL_X4 FILLER_133_1038 ();
 FILLCELL_X1 FILLER_133_1042 ();
 FILLCELL_X16 FILLER_133_1063 ();
 FILLCELL_X8 FILLER_133_1079 ();
 FILLCELL_X2 FILLER_133_1087 ();
 FILLCELL_X4 FILLER_133_1092 ();
 FILLCELL_X2 FILLER_133_1096 ();
 FILLCELL_X1 FILLER_133_1098 ();
 FILLCELL_X16 FILLER_133_1111 ();
 FILLCELL_X2 FILLER_133_1127 ();
 FILLCELL_X2 FILLER_133_1136 ();
 FILLCELL_X1 FILLER_133_1138 ();
 FILLCELL_X32 FILLER_133_1142 ();
 FILLCELL_X32 FILLER_133_1174 ();
 FILLCELL_X8 FILLER_133_1206 ();
 FILLCELL_X4 FILLER_133_1214 ();
 FILLCELL_X2 FILLER_133_1218 ();
 FILLCELL_X16 FILLER_133_1223 ();
 FILLCELL_X4 FILLER_133_1239 ();
 FILLCELL_X8 FILLER_133_1246 ();
 FILLCELL_X1 FILLER_133_1254 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X4 FILLER_134_33 ();
 FILLCELL_X2 FILLER_134_37 ();
 FILLCELL_X16 FILLER_134_46 ();
 FILLCELL_X8 FILLER_134_62 ();
 FILLCELL_X2 FILLER_134_70 ();
 FILLCELL_X16 FILLER_134_74 ();
 FILLCELL_X1 FILLER_134_104 ();
 FILLCELL_X4 FILLER_134_132 ();
 FILLCELL_X2 FILLER_134_136 ();
 FILLCELL_X4 FILLER_134_141 ();
 FILLCELL_X1 FILLER_134_145 ();
 FILLCELL_X2 FILLER_134_156 ();
 FILLCELL_X8 FILLER_134_160 ();
 FILLCELL_X4 FILLER_134_168 ();
 FILLCELL_X2 FILLER_134_172 ();
 FILLCELL_X1 FILLER_134_174 ();
 FILLCELL_X2 FILLER_134_182 ();
 FILLCELL_X1 FILLER_134_205 ();
 FILLCELL_X4 FILLER_134_209 ();
 FILLCELL_X2 FILLER_134_220 ();
 FILLCELL_X1 FILLER_134_222 ();
 FILLCELL_X1 FILLER_134_233 ();
 FILLCELL_X2 FILLER_134_260 ();
 FILLCELL_X1 FILLER_134_262 ();
 FILLCELL_X2 FILLER_134_277 ();
 FILLCELL_X2 FILLER_134_286 ();
 FILLCELL_X1 FILLER_134_288 ();
 FILLCELL_X4 FILLER_134_296 ();
 FILLCELL_X2 FILLER_134_300 ();
 FILLCELL_X8 FILLER_134_323 ();
 FILLCELL_X4 FILLER_134_331 ();
 FILLCELL_X1 FILLER_134_335 ();
 FILLCELL_X8 FILLER_134_343 ();
 FILLCELL_X1 FILLER_134_351 ();
 FILLCELL_X4 FILLER_134_359 ();
 FILLCELL_X8 FILLER_134_370 ();
 FILLCELL_X4 FILLER_134_378 ();
 FILLCELL_X1 FILLER_134_382 ();
 FILLCELL_X2 FILLER_134_410 ();
 FILLCELL_X1 FILLER_134_412 ();
 FILLCELL_X1 FILLER_134_453 ();
 FILLCELL_X1 FILLER_134_474 ();
 FILLCELL_X2 FILLER_134_494 ();
 FILLCELL_X32 FILLER_134_528 ();
 FILLCELL_X1 FILLER_134_560 ();
 FILLCELL_X8 FILLER_134_578 ();
 FILLCELL_X1 FILLER_134_596 ();
 FILLCELL_X8 FILLER_134_618 ();
 FILLCELL_X4 FILLER_134_626 ();
 FILLCELL_X1 FILLER_134_630 ();
 FILLCELL_X8 FILLER_134_632 ();
 FILLCELL_X1 FILLER_134_640 ();
 FILLCELL_X8 FILLER_134_671 ();
 FILLCELL_X2 FILLER_134_679 ();
 FILLCELL_X2 FILLER_134_708 ();
 FILLCELL_X1 FILLER_134_710 ();
 FILLCELL_X2 FILLER_134_720 ();
 FILLCELL_X1 FILLER_134_722 ();
 FILLCELL_X1 FILLER_134_730 ();
 FILLCELL_X4 FILLER_134_745 ();
 FILLCELL_X2 FILLER_134_749 ();
 FILLCELL_X8 FILLER_134_784 ();
 FILLCELL_X4 FILLER_134_792 ();
 FILLCELL_X1 FILLER_134_796 ();
 FILLCELL_X16 FILLER_134_806 ();
 FILLCELL_X8 FILLER_134_822 ();
 FILLCELL_X2 FILLER_134_830 ();
 FILLCELL_X1 FILLER_134_832 ();
 FILLCELL_X2 FILLER_134_838 ();
 FILLCELL_X8 FILLER_134_867 ();
 FILLCELL_X4 FILLER_134_875 ();
 FILLCELL_X2 FILLER_134_879 ();
 FILLCELL_X8 FILLER_134_888 ();
 FILLCELL_X2 FILLER_134_896 ();
 FILLCELL_X1 FILLER_134_905 ();
 FILLCELL_X1 FILLER_134_913 ();
 FILLCELL_X2 FILLER_134_928 ();
 FILLCELL_X1 FILLER_134_933 ();
 FILLCELL_X4 FILLER_134_954 ();
 FILLCELL_X1 FILLER_134_958 ();
 FILLCELL_X4 FILLER_134_985 ();
 FILLCELL_X16 FILLER_134_1015 ();
 FILLCELL_X8 FILLER_134_1031 ();
 FILLCELL_X4 FILLER_134_1039 ();
 FILLCELL_X2 FILLER_134_1043 ();
 FILLCELL_X2 FILLER_134_1055 ();
 FILLCELL_X4 FILLER_134_1061 ();
 FILLCELL_X4 FILLER_134_1075 ();
 FILLCELL_X4 FILLER_134_1081 ();
 FILLCELL_X2 FILLER_134_1085 ();
 FILLCELL_X1 FILLER_134_1087 ();
 FILLCELL_X2 FILLER_134_1106 ();
 FILLCELL_X4 FILLER_134_1112 ();
 FILLCELL_X2 FILLER_134_1130 ();
 FILLCELL_X1 FILLER_134_1132 ();
 FILLCELL_X4 FILLER_134_1135 ();
 FILLCELL_X32 FILLER_134_1151 ();
 FILLCELL_X32 FILLER_134_1183 ();
 FILLCELL_X16 FILLER_134_1215 ();
 FILLCELL_X8 FILLER_134_1231 ();
 FILLCELL_X1 FILLER_134_1242 ();
 FILLCELL_X2 FILLER_134_1246 ();
 FILLCELL_X1 FILLER_134_1248 ();
 FILLCELL_X2 FILLER_134_1252 ();
 FILLCELL_X1 FILLER_134_1254 ();
 FILLCELL_X16 FILLER_135_1 ();
 FILLCELL_X1 FILLER_135_17 ();
 FILLCELL_X4 FILLER_135_38 ();
 FILLCELL_X2 FILLER_135_42 ();
 FILLCELL_X1 FILLER_135_64 ();
 FILLCELL_X8 FILLER_135_79 ();
 FILLCELL_X1 FILLER_135_87 ();
 FILLCELL_X8 FILLER_135_95 ();
 FILLCELL_X2 FILLER_135_103 ();
 FILLCELL_X1 FILLER_135_105 ();
 FILLCELL_X8 FILLER_135_113 ();
 FILLCELL_X4 FILLER_135_121 ();
 FILLCELL_X2 FILLER_135_125 ();
 FILLCELL_X1 FILLER_135_127 ();
 FILLCELL_X2 FILLER_135_155 ();
 FILLCELL_X2 FILLER_135_167 ();
 FILLCELL_X4 FILLER_135_193 ();
 FILLCELL_X2 FILLER_135_204 ();
 FILLCELL_X2 FILLER_135_231 ();
 FILLCELL_X2 FILLER_135_238 ();
 FILLCELL_X8 FILLER_135_260 ();
 FILLCELL_X4 FILLER_135_268 ();
 FILLCELL_X2 FILLER_135_279 ();
 FILLCELL_X2 FILLER_135_308 ();
 FILLCELL_X1 FILLER_135_310 ();
 FILLCELL_X8 FILLER_135_318 ();
 FILLCELL_X4 FILLER_135_326 ();
 FILLCELL_X8 FILLER_135_364 ();
 FILLCELL_X2 FILLER_135_372 ();
 FILLCELL_X1 FILLER_135_374 ();
 FILLCELL_X2 FILLER_135_395 ();
 FILLCELL_X16 FILLER_135_452 ();
 FILLCELL_X8 FILLER_135_468 ();
 FILLCELL_X4 FILLER_135_476 ();
 FILLCELL_X1 FILLER_135_480 ();
 FILLCELL_X2 FILLER_135_501 ();
 FILLCELL_X8 FILLER_135_506 ();
 FILLCELL_X2 FILLER_135_521 ();
 FILLCELL_X1 FILLER_135_523 ();
 FILLCELL_X4 FILLER_135_555 ();
 FILLCELL_X4 FILLER_135_580 ();
 FILLCELL_X2 FILLER_135_584 ();
 FILLCELL_X2 FILLER_135_600 ();
 FILLCELL_X1 FILLER_135_602 ();
 FILLCELL_X4 FILLER_135_641 ();
 FILLCELL_X4 FILLER_135_673 ();
 FILLCELL_X4 FILLER_135_684 ();
 FILLCELL_X2 FILLER_135_688 ();
 FILLCELL_X1 FILLER_135_690 ();
 FILLCELL_X4 FILLER_135_705 ();
 FILLCELL_X8 FILLER_135_741 ();
 FILLCELL_X1 FILLER_135_749 ();
 FILLCELL_X8 FILLER_135_763 ();
 FILLCELL_X4 FILLER_135_771 ();
 FILLCELL_X1 FILLER_135_784 ();
 FILLCELL_X1 FILLER_135_803 ();
 FILLCELL_X2 FILLER_135_813 ();
 FILLCELL_X1 FILLER_135_815 ();
 FILLCELL_X2 FILLER_135_825 ();
 FILLCELL_X1 FILLER_135_868 ();
 FILLCELL_X1 FILLER_135_895 ();
 FILLCELL_X2 FILLER_135_903 ();
 FILLCELL_X2 FILLER_135_908 ();
 FILLCELL_X2 FILLER_135_917 ();
 FILLCELL_X1 FILLER_135_938 ();
 FILLCELL_X1 FILLER_135_943 ();
 FILLCELL_X4 FILLER_135_948 ();
 FILLCELL_X1 FILLER_135_956 ();
 FILLCELL_X1 FILLER_135_960 ();
 FILLCELL_X1 FILLER_135_965 ();
 FILLCELL_X1 FILLER_135_970 ();
 FILLCELL_X1 FILLER_135_978 ();
 FILLCELL_X1 FILLER_135_996 ();
 FILLCELL_X4 FILLER_135_1004 ();
 FILLCELL_X8 FILLER_135_1021 ();
 FILLCELL_X4 FILLER_135_1029 ();
 FILLCELL_X1 FILLER_135_1033 ();
 FILLCELL_X1 FILLER_135_1044 ();
 FILLCELL_X1 FILLER_135_1055 ();
 FILLCELL_X1 FILLER_135_1082 ();
 FILLCELL_X8 FILLER_135_1099 ();
 FILLCELL_X4 FILLER_135_1107 ();
 FILLCELL_X4 FILLER_135_1115 ();
 FILLCELL_X2 FILLER_135_1119 ();
 FILLCELL_X4 FILLER_135_1133 ();
 FILLCELL_X2 FILLER_135_1137 ();
 FILLCELL_X32 FILLER_135_1161 ();
 FILLCELL_X32 FILLER_135_1193 ();
 FILLCELL_X16 FILLER_135_1225 ();
 FILLCELL_X8 FILLER_135_1241 ();
 FILLCELL_X4 FILLER_135_1249 ();
 FILLCELL_X2 FILLER_135_1253 ();
 FILLCELL_X16 FILLER_136_1 ();
 FILLCELL_X8 FILLER_136_17 ();
 FILLCELL_X4 FILLER_136_25 ();
 FILLCELL_X8 FILLER_136_36 ();
 FILLCELL_X8 FILLER_136_51 ();
 FILLCELL_X4 FILLER_136_59 ();
 FILLCELL_X2 FILLER_136_63 ();
 FILLCELL_X4 FILLER_136_79 ();
 FILLCELL_X4 FILLER_136_110 ();
 FILLCELL_X16 FILLER_136_128 ();
 FILLCELL_X2 FILLER_136_144 ();
 FILLCELL_X1 FILLER_136_146 ();
 FILLCELL_X2 FILLER_136_154 ();
 FILLCELL_X1 FILLER_136_156 ();
 FILLCELL_X16 FILLER_136_190 ();
 FILLCELL_X8 FILLER_136_206 ();
 FILLCELL_X4 FILLER_136_214 ();
 FILLCELL_X2 FILLER_136_218 ();
 FILLCELL_X2 FILLER_136_230 ();
 FILLCELL_X1 FILLER_136_232 ();
 FILLCELL_X1 FILLER_136_240 ();
 FILLCELL_X4 FILLER_136_254 ();
 FILLCELL_X2 FILLER_136_258 ();
 FILLCELL_X1 FILLER_136_260 ();
 FILLCELL_X8 FILLER_136_281 ();
 FILLCELL_X4 FILLER_136_289 ();
 FILLCELL_X1 FILLER_136_293 ();
 FILLCELL_X4 FILLER_136_314 ();
 FILLCELL_X2 FILLER_136_318 ();
 FILLCELL_X4 FILLER_136_347 ();
 FILLCELL_X2 FILLER_136_351 ();
 FILLCELL_X1 FILLER_136_353 ();
 FILLCELL_X16 FILLER_136_361 ();
 FILLCELL_X4 FILLER_136_377 ();
 FILLCELL_X1 FILLER_136_381 ();
 FILLCELL_X1 FILLER_136_392 ();
 FILLCELL_X4 FILLER_136_416 ();
 FILLCELL_X2 FILLER_136_420 ();
 FILLCELL_X2 FILLER_136_429 ();
 FILLCELL_X8 FILLER_136_442 ();
 FILLCELL_X1 FILLER_136_450 ();
 FILLCELL_X4 FILLER_136_458 ();
 FILLCELL_X2 FILLER_136_462 ();
 FILLCELL_X1 FILLER_136_464 ();
 FILLCELL_X4 FILLER_136_476 ();
 FILLCELL_X1 FILLER_136_480 ();
 FILLCELL_X8 FILLER_136_488 ();
 FILLCELL_X1 FILLER_136_523 ();
 FILLCELL_X16 FILLER_136_531 ();
 FILLCELL_X8 FILLER_136_547 ();
 FILLCELL_X2 FILLER_136_555 ();
 FILLCELL_X1 FILLER_136_557 ();
 FILLCELL_X1 FILLER_136_590 ();
 FILLCELL_X2 FILLER_136_621 ();
 FILLCELL_X1 FILLER_136_630 ();
 FILLCELL_X2 FILLER_136_632 ();
 FILLCELL_X1 FILLER_136_634 ();
 FILLCELL_X4 FILLER_136_670 ();
 FILLCELL_X1 FILLER_136_674 ();
 FILLCELL_X8 FILLER_136_695 ();
 FILLCELL_X4 FILLER_136_703 ();
 FILLCELL_X2 FILLER_136_707 ();
 FILLCELL_X1 FILLER_136_709 ();
 FILLCELL_X8 FILLER_136_717 ();
 FILLCELL_X2 FILLER_136_725 ();
 FILLCELL_X1 FILLER_136_727 ();
 FILLCELL_X8 FILLER_136_749 ();
 FILLCELL_X4 FILLER_136_757 ();
 FILLCELL_X1 FILLER_136_761 ();
 FILLCELL_X2 FILLER_136_774 ();
 FILLCELL_X1 FILLER_136_776 ();
 FILLCELL_X4 FILLER_136_791 ();
 FILLCELL_X2 FILLER_136_795 ();
 FILLCELL_X1 FILLER_136_813 ();
 FILLCELL_X4 FILLER_136_830 ();
 FILLCELL_X2 FILLER_136_871 ();
 FILLCELL_X1 FILLER_136_880 ();
 FILLCELL_X4 FILLER_136_891 ();
 FILLCELL_X2 FILLER_136_915 ();
 FILLCELL_X4 FILLER_136_944 ();
 FILLCELL_X1 FILLER_136_948 ();
 FILLCELL_X1 FILLER_136_975 ();
 FILLCELL_X2 FILLER_136_1003 ();
 FILLCELL_X2 FILLER_136_1009 ();
 FILLCELL_X1 FILLER_136_1011 ();
 FILLCELL_X4 FILLER_136_1021 ();
 FILLCELL_X1 FILLER_136_1025 ();
 FILLCELL_X2 FILLER_136_1036 ();
 FILLCELL_X1 FILLER_136_1068 ();
 FILLCELL_X1 FILLER_136_1071 ();
 FILLCELL_X1 FILLER_136_1074 ();
 FILLCELL_X4 FILLER_136_1087 ();
 FILLCELL_X1 FILLER_136_1091 ();
 FILLCELL_X4 FILLER_136_1124 ();
 FILLCELL_X2 FILLER_136_1128 ();
 FILLCELL_X4 FILLER_136_1132 ();
 FILLCELL_X2 FILLER_136_1138 ();
 FILLCELL_X1 FILLER_136_1140 ();
 FILLCELL_X8 FILLER_136_1151 ();
 FILLCELL_X2 FILLER_136_1159 ();
 FILLCELL_X32 FILLER_136_1173 ();
 FILLCELL_X32 FILLER_136_1205 ();
 FILLCELL_X16 FILLER_136_1237 ();
 FILLCELL_X2 FILLER_136_1253 ();
 FILLCELL_X16 FILLER_137_1 ();
 FILLCELL_X1 FILLER_137_17 ();
 FILLCELL_X1 FILLER_137_38 ();
 FILLCELL_X2 FILLER_137_66 ();
 FILLCELL_X4 FILLER_137_75 ();
 FILLCELL_X2 FILLER_137_79 ();
 FILLCELL_X4 FILLER_137_101 ();
 FILLCELL_X1 FILLER_137_105 ();
 FILLCELL_X8 FILLER_137_113 ();
 FILLCELL_X1 FILLER_137_121 ();
 FILLCELL_X4 FILLER_137_129 ();
 FILLCELL_X2 FILLER_137_133 ();
 FILLCELL_X8 FILLER_137_175 ();
 FILLCELL_X2 FILLER_137_183 ();
 FILLCELL_X2 FILLER_137_192 ();
 FILLCELL_X2 FILLER_137_221 ();
 FILLCELL_X1 FILLER_137_223 ();
 FILLCELL_X4 FILLER_137_244 ();
 FILLCELL_X2 FILLER_137_248 ();
 FILLCELL_X2 FILLER_137_270 ();
 FILLCELL_X1 FILLER_137_272 ();
 FILLCELL_X2 FILLER_137_280 ();
 FILLCELL_X2 FILLER_137_286 ();
 FILLCELL_X1 FILLER_137_288 ();
 FILLCELL_X4 FILLER_137_293 ();
 FILLCELL_X1 FILLER_137_321 ();
 FILLCELL_X2 FILLER_137_349 ();
 FILLCELL_X1 FILLER_137_351 ();
 FILLCELL_X4 FILLER_137_366 ();
 FILLCELL_X2 FILLER_137_370 ();
 FILLCELL_X1 FILLER_137_372 ();
 FILLCELL_X2 FILLER_137_405 ();
 FILLCELL_X2 FILLER_137_416 ();
 FILLCELL_X4 FILLER_137_438 ();
 FILLCELL_X1 FILLER_137_442 ();
 FILLCELL_X4 FILLER_137_470 ();
 FILLCELL_X1 FILLER_137_474 ();
 FILLCELL_X16 FILLER_137_493 ();
 FILLCELL_X8 FILLER_137_509 ();
 FILLCELL_X4 FILLER_137_517 ();
 FILLCELL_X1 FILLER_137_521 ();
 FILLCELL_X4 FILLER_137_531 ();
 FILLCELL_X2 FILLER_137_542 ();
 FILLCELL_X1 FILLER_137_544 ();
 FILLCELL_X4 FILLER_137_572 ();
 FILLCELL_X1 FILLER_137_576 ();
 FILLCELL_X4 FILLER_137_590 ();
 FILLCELL_X1 FILLER_137_594 ();
 FILLCELL_X8 FILLER_137_602 ();
 FILLCELL_X4 FILLER_137_610 ();
 FILLCELL_X2 FILLER_137_614 ();
 FILLCELL_X1 FILLER_137_616 ();
 FILLCELL_X2 FILLER_137_645 ();
 FILLCELL_X1 FILLER_137_647 ();
 FILLCELL_X8 FILLER_137_672 ();
 FILLCELL_X2 FILLER_137_680 ();
 FILLCELL_X1 FILLER_137_682 ();
 FILLCELL_X16 FILLER_137_695 ();
 FILLCELL_X4 FILLER_137_711 ();
 FILLCELL_X32 FILLER_137_722 ();
 FILLCELL_X2 FILLER_137_754 ();
 FILLCELL_X1 FILLER_137_756 ();
 FILLCELL_X1 FILLER_137_799 ();
 FILLCELL_X2 FILLER_137_826 ();
 FILLCELL_X1 FILLER_137_828 ();
 FILLCELL_X4 FILLER_137_836 ();
 FILLCELL_X2 FILLER_137_840 ();
 FILLCELL_X1 FILLER_137_842 ();
 FILLCELL_X2 FILLER_137_882 ();
 FILLCELL_X4 FILLER_137_913 ();
 FILLCELL_X1 FILLER_137_926 ();
 FILLCELL_X4 FILLER_137_940 ();
 FILLCELL_X2 FILLER_137_944 ();
 FILLCELL_X4 FILLER_137_950 ();
 FILLCELL_X2 FILLER_137_954 ();
 FILLCELL_X1 FILLER_137_956 ();
 FILLCELL_X2 FILLER_137_996 ();
 FILLCELL_X1 FILLER_137_998 ();
 FILLCELL_X1 FILLER_137_1013 ();
 FILLCELL_X1 FILLER_137_1017 ();
 FILLCELL_X2 FILLER_137_1036 ();
 FILLCELL_X4 FILLER_137_1050 ();
 FILLCELL_X2 FILLER_137_1054 ();
 FILLCELL_X2 FILLER_137_1072 ();
 FILLCELL_X1 FILLER_137_1074 ();
 FILLCELL_X4 FILLER_137_1085 ();
 FILLCELL_X2 FILLER_137_1089 ();
 FILLCELL_X2 FILLER_137_1101 ();
 FILLCELL_X2 FILLER_137_1145 ();
 FILLCELL_X1 FILLER_137_1160 ();
 FILLCELL_X32 FILLER_137_1174 ();
 FILLCELL_X32 FILLER_137_1206 ();
 FILLCELL_X16 FILLER_137_1238 ();
 FILLCELL_X1 FILLER_137_1254 ();
 FILLCELL_X16 FILLER_138_1 ();
 FILLCELL_X8 FILLER_138_17 ();
 FILLCELL_X4 FILLER_138_25 ();
 FILLCELL_X2 FILLER_138_36 ();
 FILLCELL_X4 FILLER_138_45 ();
 FILLCELL_X1 FILLER_138_49 ();
 FILLCELL_X16 FILLER_138_62 ();
 FILLCELL_X4 FILLER_138_78 ();
 FILLCELL_X2 FILLER_138_116 ();
 FILLCELL_X8 FILLER_138_125 ();
 FILLCELL_X4 FILLER_138_133 ();
 FILLCELL_X2 FILLER_138_137 ();
 FILLCELL_X1 FILLER_138_139 ();
 FILLCELL_X4 FILLER_138_143 ();
 FILLCELL_X1 FILLER_138_147 ();
 FILLCELL_X1 FILLER_138_153 ();
 FILLCELL_X8 FILLER_138_168 ();
 FILLCELL_X1 FILLER_138_176 ();
 FILLCELL_X1 FILLER_138_210 ();
 FILLCELL_X1 FILLER_138_218 ();
 FILLCELL_X1 FILLER_138_230 ();
 FILLCELL_X8 FILLER_138_246 ();
 FILLCELL_X4 FILLER_138_254 ();
 FILLCELL_X1 FILLER_138_258 ();
 FILLCELL_X8 FILLER_138_273 ();
 FILLCELL_X4 FILLER_138_305 ();
 FILLCELL_X4 FILLER_138_328 ();
 FILLCELL_X1 FILLER_138_332 ();
 FILLCELL_X4 FILLER_138_380 ();
 FILLCELL_X1 FILLER_138_384 ();
 FILLCELL_X1 FILLER_138_413 ();
 FILLCELL_X1 FILLER_138_421 ();
 FILLCELL_X16 FILLER_138_433 ();
 FILLCELL_X8 FILLER_138_449 ();
 FILLCELL_X2 FILLER_138_457 ();
 FILLCELL_X1 FILLER_138_459 ();
 FILLCELL_X2 FILLER_138_467 ();
 FILLCELL_X16 FILLER_138_487 ();
 FILLCELL_X1 FILLER_138_503 ();
 FILLCELL_X8 FILLER_138_511 ();
 FILLCELL_X2 FILLER_138_519 ();
 FILLCELL_X2 FILLER_138_546 ();
 FILLCELL_X1 FILLER_138_548 ();
 FILLCELL_X4 FILLER_138_556 ();
 FILLCELL_X1 FILLER_138_560 ();
 FILLCELL_X4 FILLER_138_581 ();
 FILLCELL_X1 FILLER_138_585 ();
 FILLCELL_X2 FILLER_138_600 ();
 FILLCELL_X1 FILLER_138_602 ();
 FILLCELL_X1 FILLER_138_606 ();
 FILLCELL_X2 FILLER_138_632 ();
 FILLCELL_X1 FILLER_138_634 ();
 FILLCELL_X2 FILLER_138_656 ();
 FILLCELL_X1 FILLER_138_672 ();
 FILLCELL_X2 FILLER_138_747 ();
 FILLCELL_X1 FILLER_138_758 ();
 FILLCELL_X4 FILLER_138_780 ();
 FILLCELL_X2 FILLER_138_784 ();
 FILLCELL_X1 FILLER_138_793 ();
 FILLCELL_X1 FILLER_138_811 ();
 FILLCELL_X2 FILLER_138_821 ();
 FILLCELL_X4 FILLER_138_837 ();
 FILLCELL_X1 FILLER_138_841 ();
 FILLCELL_X8 FILLER_138_847 ();
 FILLCELL_X2 FILLER_138_855 ();
 FILLCELL_X1 FILLER_138_857 ();
 FILLCELL_X8 FILLER_138_871 ();
 FILLCELL_X1 FILLER_138_879 ();
 FILLCELL_X2 FILLER_138_890 ();
 FILLCELL_X1 FILLER_138_892 ();
 FILLCELL_X1 FILLER_138_898 ();
 FILLCELL_X1 FILLER_138_913 ();
 FILLCELL_X1 FILLER_138_921 ();
 FILLCELL_X4 FILLER_138_939 ();
 FILLCELL_X2 FILLER_138_952 ();
 FILLCELL_X1 FILLER_138_954 ();
 FILLCELL_X2 FILLER_138_960 ();
 FILLCELL_X1 FILLER_138_962 ();
 FILLCELL_X1 FILLER_138_967 ();
 FILLCELL_X1 FILLER_138_976 ();
 FILLCELL_X4 FILLER_138_985 ();
 FILLCELL_X8 FILLER_138_993 ();
 FILLCELL_X2 FILLER_138_1001 ();
 FILLCELL_X1 FILLER_138_1003 ();
 FILLCELL_X8 FILLER_138_1006 ();
 FILLCELL_X1 FILLER_138_1014 ();
 FILLCELL_X8 FILLER_138_1017 ();
 FILLCELL_X2 FILLER_138_1025 ();
 FILLCELL_X1 FILLER_138_1027 ();
 FILLCELL_X2 FILLER_138_1041 ();
 FILLCELL_X1 FILLER_138_1062 ();
 FILLCELL_X4 FILLER_138_1065 ();
 FILLCELL_X2 FILLER_138_1069 ();
 FILLCELL_X8 FILLER_138_1081 ();
 FILLCELL_X2 FILLER_138_1089 ();
 FILLCELL_X4 FILLER_138_1093 ();
 FILLCELL_X1 FILLER_138_1097 ();
 FILLCELL_X16 FILLER_138_1108 ();
 FILLCELL_X8 FILLER_138_1124 ();
 FILLCELL_X2 FILLER_138_1132 ();
 FILLCELL_X1 FILLER_138_1134 ();
 FILLCELL_X8 FILLER_138_1149 ();
 FILLCELL_X4 FILLER_138_1157 ();
 FILLCELL_X2 FILLER_138_1161 ();
 FILLCELL_X32 FILLER_138_1185 ();
 FILLCELL_X32 FILLER_138_1217 ();
 FILLCELL_X4 FILLER_138_1249 ();
 FILLCELL_X2 FILLER_138_1253 ();
 FILLCELL_X16 FILLER_139_1 ();
 FILLCELL_X8 FILLER_139_17 ();
 FILLCELL_X2 FILLER_139_25 ();
 FILLCELL_X4 FILLER_139_47 ();
 FILLCELL_X4 FILLER_139_85 ();
 FILLCELL_X4 FILLER_139_96 ();
 FILLCELL_X1 FILLER_139_100 ();
 FILLCELL_X4 FILLER_139_148 ();
 FILLCELL_X4 FILLER_139_207 ();
 FILLCELL_X1 FILLER_139_211 ();
 FILLCELL_X16 FILLER_139_243 ();
 FILLCELL_X1 FILLER_139_259 ();
 FILLCELL_X16 FILLER_139_287 ();
 FILLCELL_X2 FILLER_139_303 ();
 FILLCELL_X1 FILLER_139_305 ();
 FILLCELL_X32 FILLER_139_320 ();
 FILLCELL_X1 FILLER_139_352 ();
 FILLCELL_X8 FILLER_139_360 ();
 FILLCELL_X2 FILLER_139_368 ();
 FILLCELL_X16 FILLER_139_377 ();
 FILLCELL_X1 FILLER_139_393 ();
 FILLCELL_X1 FILLER_139_401 ();
 FILLCELL_X8 FILLER_139_409 ();
 FILLCELL_X2 FILLER_139_417 ();
 FILLCELL_X1 FILLER_139_419 ();
 FILLCELL_X2 FILLER_139_468 ();
 FILLCELL_X4 FILLER_139_477 ();
 FILLCELL_X4 FILLER_139_488 ();
 FILLCELL_X2 FILLER_139_492 ();
 FILLCELL_X4 FILLER_139_528 ();
 FILLCELL_X2 FILLER_139_546 ();
 FILLCELL_X1 FILLER_139_548 ();
 FILLCELL_X2 FILLER_139_569 ();
 FILLCELL_X1 FILLER_139_571 ();
 FILLCELL_X16 FILLER_139_579 ();
 FILLCELL_X1 FILLER_139_615 ();
 FILLCELL_X1 FILLER_139_630 ();
 FILLCELL_X1 FILLER_139_634 ();
 FILLCELL_X1 FILLER_139_642 ();
 FILLCELL_X1 FILLER_139_646 ();
 FILLCELL_X2 FILLER_139_661 ();
 FILLCELL_X2 FILLER_139_676 ();
 FILLCELL_X1 FILLER_139_678 ();
 FILLCELL_X2 FILLER_139_699 ();
 FILLCELL_X1 FILLER_139_701 ();
 FILLCELL_X2 FILLER_139_709 ();
 FILLCELL_X1 FILLER_139_711 ();
 FILLCELL_X4 FILLER_139_726 ();
 FILLCELL_X2 FILLER_139_730 ();
 FILLCELL_X1 FILLER_139_732 ();
 FILLCELL_X1 FILLER_139_740 ();
 FILLCELL_X8 FILLER_139_778 ();
 FILLCELL_X4 FILLER_139_786 ();
 FILLCELL_X1 FILLER_139_790 ();
 FILLCELL_X2 FILLER_139_798 ();
 FILLCELL_X1 FILLER_139_800 ();
 FILLCELL_X4 FILLER_139_804 ();
 FILLCELL_X2 FILLER_139_808 ();
 FILLCELL_X1 FILLER_139_810 ();
 FILLCELL_X2 FILLER_139_820 ();
 FILLCELL_X1 FILLER_139_822 ();
 FILLCELL_X4 FILLER_139_832 ();
 FILLCELL_X2 FILLER_139_836 ();
 FILLCELL_X1 FILLER_139_838 ();
 FILLCELL_X2 FILLER_139_849 ();
 FILLCELL_X1 FILLER_139_855 ();
 FILLCELL_X8 FILLER_139_860 ();
 FILLCELL_X4 FILLER_139_868 ();
 FILLCELL_X1 FILLER_139_872 ();
 FILLCELL_X16 FILLER_139_887 ();
 FILLCELL_X2 FILLER_139_910 ();
 FILLCELL_X1 FILLER_139_912 ();
 FILLCELL_X8 FILLER_139_916 ();
 FILLCELL_X1 FILLER_139_924 ();
 FILLCELL_X16 FILLER_139_940 ();
 FILLCELL_X4 FILLER_139_956 ();
 FILLCELL_X2 FILLER_139_960 ();
 FILLCELL_X1 FILLER_139_962 ();
 FILLCELL_X2 FILLER_139_967 ();
 FILLCELL_X4 FILLER_139_978 ();
 FILLCELL_X2 FILLER_139_1001 ();
 FILLCELL_X1 FILLER_139_1005 ();
 FILLCELL_X8 FILLER_139_1031 ();
 FILLCELL_X2 FILLER_139_1039 ();
 FILLCELL_X4 FILLER_139_1059 ();
 FILLCELL_X2 FILLER_139_1063 ();
 FILLCELL_X1 FILLER_139_1065 ();
 FILLCELL_X4 FILLER_139_1071 ();
 FILLCELL_X2 FILLER_139_1075 ();
 FILLCELL_X1 FILLER_139_1077 ();
 FILLCELL_X8 FILLER_139_1080 ();
 FILLCELL_X1 FILLER_139_1088 ();
 FILLCELL_X2 FILLER_139_1091 ();
 FILLCELL_X1 FILLER_139_1120 ();
 FILLCELL_X4 FILLER_139_1123 ();
 FILLCELL_X2 FILLER_139_1127 ();
 FILLCELL_X1 FILLER_139_1129 ();
 FILLCELL_X1 FILLER_139_1142 ();
 FILLCELL_X4 FILLER_139_1159 ();
 FILLCELL_X1 FILLER_139_1167 ();
 FILLCELL_X2 FILLER_139_1171 ();
 FILLCELL_X32 FILLER_139_1180 ();
 FILLCELL_X32 FILLER_139_1212 ();
 FILLCELL_X8 FILLER_139_1244 ();
 FILLCELL_X2 FILLER_139_1252 ();
 FILLCELL_X1 FILLER_139_1254 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X4 FILLER_140_33 ();
 FILLCELL_X2 FILLER_140_37 ();
 FILLCELL_X1 FILLER_140_39 ();
 FILLCELL_X8 FILLER_140_47 ();
 FILLCELL_X2 FILLER_140_62 ();
 FILLCELL_X2 FILLER_140_71 ();
 FILLCELL_X1 FILLER_140_73 ();
 FILLCELL_X2 FILLER_140_81 ();
 FILLCELL_X1 FILLER_140_83 ();
 FILLCELL_X16 FILLER_140_91 ();
 FILLCELL_X8 FILLER_140_114 ();
 FILLCELL_X4 FILLER_140_122 ();
 FILLCELL_X1 FILLER_140_126 ();
 FILLCELL_X4 FILLER_140_134 ();
 FILLCELL_X2 FILLER_140_138 ();
 FILLCELL_X8 FILLER_140_167 ();
 FILLCELL_X4 FILLER_140_175 ();
 FILLCELL_X4 FILLER_140_193 ();
 FILLCELL_X2 FILLER_140_197 ();
 FILLCELL_X1 FILLER_140_199 ();
 FILLCELL_X16 FILLER_140_220 ();
 FILLCELL_X2 FILLER_140_236 ();
 FILLCELL_X8 FILLER_140_243 ();
 FILLCELL_X2 FILLER_140_251 ();
 FILLCELL_X1 FILLER_140_253 ();
 FILLCELL_X4 FILLER_140_308 ();
 FILLCELL_X2 FILLER_140_312 ();
 FILLCELL_X4 FILLER_140_321 ();
 FILLCELL_X8 FILLER_140_359 ();
 FILLCELL_X8 FILLER_140_387 ();
 FILLCELL_X4 FILLER_140_395 ();
 FILLCELL_X1 FILLER_140_399 ();
 FILLCELL_X8 FILLER_140_407 ();
 FILLCELL_X2 FILLER_140_415 ();
 FILLCELL_X1 FILLER_140_417 ();
 FILLCELL_X4 FILLER_140_445 ();
 FILLCELL_X2 FILLER_140_449 ();
 FILLCELL_X1 FILLER_140_451 ();
 FILLCELL_X4 FILLER_140_459 ();
 FILLCELL_X4 FILLER_140_466 ();
 FILLCELL_X16 FILLER_140_507 ();
 FILLCELL_X4 FILLER_140_523 ();
 FILLCELL_X2 FILLER_140_527 ();
 FILLCELL_X1 FILLER_140_543 ();
 FILLCELL_X16 FILLER_140_571 ();
 FILLCELL_X8 FILLER_140_587 ();
 FILLCELL_X8 FILLER_140_602 ();
 FILLCELL_X2 FILLER_140_610 ();
 FILLCELL_X1 FILLER_140_619 ();
 FILLCELL_X4 FILLER_140_627 ();
 FILLCELL_X8 FILLER_140_632 ();
 FILLCELL_X2 FILLER_140_640 ();
 FILLCELL_X1 FILLER_140_642 ();
 FILLCELL_X8 FILLER_140_650 ();
 FILLCELL_X4 FILLER_140_658 ();
 FILLCELL_X1 FILLER_140_662 ();
 FILLCELL_X16 FILLER_140_666 ();
 FILLCELL_X8 FILLER_140_682 ();
 FILLCELL_X4 FILLER_140_690 ();
 FILLCELL_X2 FILLER_140_694 ();
 FILLCELL_X2 FILLER_140_716 ();
 FILLCELL_X8 FILLER_140_738 ();
 FILLCELL_X4 FILLER_140_746 ();
 FILLCELL_X2 FILLER_140_750 ();
 FILLCELL_X2 FILLER_140_768 ();
 FILLCELL_X4 FILLER_140_777 ();
 FILLCELL_X2 FILLER_140_781 ();
 FILLCELL_X1 FILLER_140_783 ();
 FILLCELL_X4 FILLER_140_791 ();
 FILLCELL_X1 FILLER_140_795 ();
 FILLCELL_X1 FILLER_140_820 ();
 FILLCELL_X4 FILLER_140_824 ();
 FILLCELL_X1 FILLER_140_828 ();
 FILLCELL_X2 FILLER_140_836 ();
 FILLCELL_X1 FILLER_140_838 ();
 FILLCELL_X2 FILLER_140_881 ();
 FILLCELL_X1 FILLER_140_883 ();
 FILLCELL_X4 FILLER_140_909 ();
 FILLCELL_X2 FILLER_140_916 ();
 FILLCELL_X2 FILLER_140_934 ();
 FILLCELL_X8 FILLER_140_953 ();
 FILLCELL_X4 FILLER_140_961 ();
 FILLCELL_X2 FILLER_140_974 ();
 FILLCELL_X1 FILLER_140_1018 ();
 FILLCELL_X2 FILLER_140_1041 ();
 FILLCELL_X1 FILLER_140_1043 ();
 FILLCELL_X1 FILLER_140_1047 ();
 FILLCELL_X1 FILLER_140_1054 ();
 FILLCELL_X1 FILLER_140_1090 ();
 FILLCELL_X2 FILLER_140_1095 ();
 FILLCELL_X1 FILLER_140_1097 ();
 FILLCELL_X1 FILLER_140_1129 ();
 FILLCELL_X2 FILLER_140_1132 ();
 FILLCELL_X8 FILLER_140_1150 ();
 FILLCELL_X4 FILLER_140_1158 ();
 FILLCELL_X1 FILLER_140_1162 ();
 FILLCELL_X1 FILLER_140_1168 ();
 FILLCELL_X32 FILLER_140_1185 ();
 FILLCELL_X32 FILLER_140_1217 ();
 FILLCELL_X4 FILLER_140_1249 ();
 FILLCELL_X2 FILLER_140_1253 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X2 FILLER_141_33 ();
 FILLCELL_X4 FILLER_141_89 ();
 FILLCELL_X1 FILLER_141_93 ();
 FILLCELL_X1 FILLER_141_121 ();
 FILLCELL_X4 FILLER_141_136 ();
 FILLCELL_X2 FILLER_141_140 ();
 FILLCELL_X1 FILLER_141_142 ();
 FILLCELL_X2 FILLER_141_150 ();
 FILLCELL_X1 FILLER_141_152 ();
 FILLCELL_X16 FILLER_141_194 ();
 FILLCELL_X8 FILLER_141_210 ();
 FILLCELL_X4 FILLER_141_218 ();
 FILLCELL_X2 FILLER_141_222 ();
 FILLCELL_X1 FILLER_141_224 ();
 FILLCELL_X8 FILLER_141_232 ();
 FILLCELL_X2 FILLER_141_240 ();
 FILLCELL_X1 FILLER_141_242 ();
 FILLCELL_X32 FILLER_141_250 ();
 FILLCELL_X2 FILLER_141_282 ();
 FILLCELL_X2 FILLER_141_291 ();
 FILLCELL_X1 FILLER_141_320 ();
 FILLCELL_X2 FILLER_141_341 ();
 FILLCELL_X1 FILLER_141_343 ();
 FILLCELL_X2 FILLER_141_358 ();
 FILLCELL_X1 FILLER_141_360 ();
 FILLCELL_X2 FILLER_141_368 ();
 FILLCELL_X2 FILLER_141_377 ();
 FILLCELL_X1 FILLER_141_379 ();
 FILLCELL_X32 FILLER_141_400 ();
 FILLCELL_X2 FILLER_141_432 ();
 FILLCELL_X1 FILLER_141_434 ();
 FILLCELL_X2 FILLER_141_479 ();
 FILLCELL_X4 FILLER_141_488 ();
 FILLCELL_X8 FILLER_141_526 ();
 FILLCELL_X2 FILLER_141_545 ();
 FILLCELL_X1 FILLER_141_547 ();
 FILLCELL_X32 FILLER_141_555 ();
 FILLCELL_X32 FILLER_141_587 ();
 FILLCELL_X32 FILLER_141_619 ();
 FILLCELL_X32 FILLER_141_651 ();
 FILLCELL_X32 FILLER_141_683 ();
 FILLCELL_X2 FILLER_141_715 ();
 FILLCELL_X1 FILLER_141_717 ();
 FILLCELL_X2 FILLER_141_734 ();
 FILLCELL_X1 FILLER_141_736 ();
 FILLCELL_X1 FILLER_141_759 ();
 FILLCELL_X8 FILLER_141_772 ();
 FILLCELL_X1 FILLER_141_780 ();
 FILLCELL_X1 FILLER_141_810 ();
 FILLCELL_X8 FILLER_141_818 ();
 FILLCELL_X2 FILLER_141_826 ();
 FILLCELL_X1 FILLER_141_828 ();
 FILLCELL_X4 FILLER_141_858 ();
 FILLCELL_X2 FILLER_141_862 ();
 FILLCELL_X1 FILLER_141_871 ();
 FILLCELL_X8 FILLER_141_879 ();
 FILLCELL_X1 FILLER_141_887 ();
 FILLCELL_X2 FILLER_141_895 ();
 FILLCELL_X1 FILLER_141_897 ();
 FILLCELL_X8 FILLER_141_918 ();
 FILLCELL_X2 FILLER_141_926 ();
 FILLCELL_X1 FILLER_141_970 ();
 FILLCELL_X8 FILLER_141_978 ();
 FILLCELL_X4 FILLER_141_986 ();
 FILLCELL_X4 FILLER_141_1000 ();
 FILLCELL_X2 FILLER_141_1004 ();
 FILLCELL_X1 FILLER_141_1006 ();
 FILLCELL_X2 FILLER_141_1059 ();
 FILLCELL_X2 FILLER_141_1064 ();
 FILLCELL_X4 FILLER_141_1069 ();
 FILLCELL_X2 FILLER_141_1073 ();
 FILLCELL_X2 FILLER_141_1094 ();
 FILLCELL_X1 FILLER_141_1096 ();
 FILLCELL_X16 FILLER_141_1110 ();
 FILLCELL_X2 FILLER_141_1126 ();
 FILLCELL_X1 FILLER_141_1128 ();
 FILLCELL_X4 FILLER_141_1133 ();
 FILLCELL_X2 FILLER_141_1137 ();
 FILLCELL_X1 FILLER_141_1139 ();
 FILLCELL_X4 FILLER_141_1150 ();
 FILLCELL_X1 FILLER_141_1164 ();
 FILLCELL_X2 FILLER_141_1169 ();
 FILLCELL_X1 FILLER_141_1171 ();
 FILLCELL_X32 FILLER_141_1181 ();
 FILLCELL_X32 FILLER_141_1213 ();
 FILLCELL_X8 FILLER_141_1245 ();
 FILLCELL_X2 FILLER_141_1253 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X4 FILLER_142_65 ();
 FILLCELL_X2 FILLER_142_69 ();
 FILLCELL_X1 FILLER_142_71 ();
 FILLCELL_X2 FILLER_142_79 ();
 FILLCELL_X1 FILLER_142_101 ();
 FILLCELL_X4 FILLER_142_137 ();
 FILLCELL_X2 FILLER_142_141 ();
 FILLCELL_X1 FILLER_142_143 ();
 FILLCELL_X2 FILLER_142_151 ();
 FILLCELL_X8 FILLER_142_167 ();
 FILLCELL_X4 FILLER_142_175 ();
 FILLCELL_X1 FILLER_142_179 ();
 FILLCELL_X1 FILLER_142_242 ();
 FILLCELL_X8 FILLER_142_263 ();
 FILLCELL_X1 FILLER_142_271 ();
 FILLCELL_X8 FILLER_142_292 ();
 FILLCELL_X4 FILLER_142_300 ();
 FILLCELL_X8 FILLER_142_311 ();
 FILLCELL_X4 FILLER_142_319 ();
 FILLCELL_X8 FILLER_142_340 ();
 FILLCELL_X8 FILLER_142_375 ();
 FILLCELL_X2 FILLER_142_383 ();
 FILLCELL_X1 FILLER_142_385 ();
 FILLCELL_X4 FILLER_142_400 ();
 FILLCELL_X16 FILLER_142_431 ();
 FILLCELL_X4 FILLER_142_447 ();
 FILLCELL_X2 FILLER_142_451 ();
 FILLCELL_X1 FILLER_142_453 ();
 FILLCELL_X1 FILLER_142_475 ();
 FILLCELL_X1 FILLER_142_479 ();
 FILLCELL_X2 FILLER_142_494 ();
 FILLCELL_X1 FILLER_142_496 ();
 FILLCELL_X4 FILLER_142_529 ();
 FILLCELL_X1 FILLER_142_533 ();
 FILLCELL_X32 FILLER_142_558 ();
 FILLCELL_X32 FILLER_142_590 ();
 FILLCELL_X8 FILLER_142_622 ();
 FILLCELL_X1 FILLER_142_630 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X8 FILLER_142_728 ();
 FILLCELL_X2 FILLER_142_736 ();
 FILLCELL_X1 FILLER_142_738 ();
 FILLCELL_X2 FILLER_142_752 ();
 FILLCELL_X1 FILLER_142_754 ();
 FILLCELL_X2 FILLER_142_762 ();
 FILLCELL_X8 FILLER_142_784 ();
 FILLCELL_X2 FILLER_142_792 ();
 FILLCELL_X1 FILLER_142_794 ();
 FILLCELL_X1 FILLER_142_801 ();
 FILLCELL_X1 FILLER_142_814 ();
 FILLCELL_X4 FILLER_142_819 ();
 FILLCELL_X1 FILLER_142_823 ();
 FILLCELL_X2 FILLER_142_841 ();
 FILLCELL_X1 FILLER_142_843 ();
 FILLCELL_X1 FILLER_142_848 ();
 FILLCELL_X4 FILLER_142_872 ();
 FILLCELL_X1 FILLER_142_876 ();
 FILLCELL_X1 FILLER_142_894 ();
 FILLCELL_X1 FILLER_142_899 ();
 FILLCELL_X2 FILLER_142_907 ();
 FILLCELL_X1 FILLER_142_913 ();
 FILLCELL_X1 FILLER_142_918 ();
 FILLCELL_X1 FILLER_142_927 ();
 FILLCELL_X4 FILLER_142_932 ();
 FILLCELL_X2 FILLER_142_936 ();
 FILLCELL_X4 FILLER_142_948 ();
 FILLCELL_X2 FILLER_142_952 ();
 FILLCELL_X1 FILLER_142_954 ();
 FILLCELL_X4 FILLER_142_958 ();
 FILLCELL_X8 FILLER_142_973 ();
 FILLCELL_X4 FILLER_142_981 ();
 FILLCELL_X4 FILLER_142_995 ();
 FILLCELL_X2 FILLER_142_1013 ();
 FILLCELL_X2 FILLER_142_1018 ();
 FILLCELL_X1 FILLER_142_1020 ();
 FILLCELL_X4 FILLER_142_1043 ();
 FILLCELL_X1 FILLER_142_1047 ();
 FILLCELL_X8 FILLER_142_1051 ();
 FILLCELL_X2 FILLER_142_1084 ();
 FILLCELL_X2 FILLER_142_1089 ();
 FILLCELL_X4 FILLER_142_1093 ();
 FILLCELL_X2 FILLER_142_1097 ();
 FILLCELL_X1 FILLER_142_1099 ();
 FILLCELL_X4 FILLER_142_1110 ();
 FILLCELL_X2 FILLER_142_1114 ();
 FILLCELL_X16 FILLER_142_1146 ();
 FILLCELL_X4 FILLER_142_1166 ();
 FILLCELL_X1 FILLER_142_1170 ();
 FILLCELL_X32 FILLER_142_1192 ();
 FILLCELL_X16 FILLER_142_1224 ();
 FILLCELL_X8 FILLER_142_1240 ();
 FILLCELL_X4 FILLER_142_1248 ();
 FILLCELL_X2 FILLER_142_1252 ();
 FILLCELL_X1 FILLER_142_1254 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X16 FILLER_143_33 ();
 FILLCELL_X8 FILLER_143_49 ();
 FILLCELL_X4 FILLER_143_57 ();
 FILLCELL_X2 FILLER_143_61 ();
 FILLCELL_X1 FILLER_143_63 ();
 FILLCELL_X8 FILLER_143_84 ();
 FILLCELL_X2 FILLER_143_92 ();
 FILLCELL_X1 FILLER_143_94 ();
 FILLCELL_X1 FILLER_143_102 ();
 FILLCELL_X4 FILLER_143_123 ();
 FILLCELL_X1 FILLER_143_134 ();
 FILLCELL_X4 FILLER_143_176 ();
 FILLCELL_X1 FILLER_143_180 ();
 FILLCELL_X2 FILLER_143_188 ();
 FILLCELL_X2 FILLER_143_197 ();
 FILLCELL_X1 FILLER_143_199 ();
 FILLCELL_X2 FILLER_143_220 ();
 FILLCELL_X1 FILLER_143_222 ();
 FILLCELL_X2 FILLER_143_230 ();
 FILLCELL_X8 FILLER_143_259 ();
 FILLCELL_X2 FILLER_143_267 ();
 FILLCELL_X1 FILLER_143_269 ();
 FILLCELL_X2 FILLER_143_290 ();
 FILLCELL_X1 FILLER_143_299 ();
 FILLCELL_X4 FILLER_143_307 ();
 FILLCELL_X2 FILLER_143_311 ();
 FILLCELL_X1 FILLER_143_313 ();
 FILLCELL_X2 FILLER_143_334 ();
 FILLCELL_X4 FILLER_143_363 ();
 FILLCELL_X2 FILLER_143_367 ();
 FILLCELL_X1 FILLER_143_369 ();
 FILLCELL_X1 FILLER_143_411 ();
 FILLCELL_X2 FILLER_143_433 ();
 FILLCELL_X1 FILLER_143_435 ();
 FILLCELL_X8 FILLER_143_456 ();
 FILLCELL_X1 FILLER_143_467 ();
 FILLCELL_X4 FILLER_143_519 ();
 FILLCELL_X1 FILLER_143_523 ();
 FILLCELL_X32 FILLER_143_578 ();
 FILLCELL_X32 FILLER_143_610 ();
 FILLCELL_X32 FILLER_143_642 ();
 FILLCELL_X16 FILLER_143_674 ();
 FILLCELL_X8 FILLER_143_690 ();
 FILLCELL_X4 FILLER_143_698 ();
 FILLCELL_X2 FILLER_143_702 ();
 FILLCELL_X1 FILLER_143_704 ();
 FILLCELL_X1 FILLER_143_753 ();
 FILLCELL_X2 FILLER_143_786 ();
 FILLCELL_X2 FILLER_143_792 ();
 FILLCELL_X1 FILLER_143_794 ();
 FILLCELL_X8 FILLER_143_801 ();
 FILLCELL_X1 FILLER_143_809 ();
 FILLCELL_X4 FILLER_143_814 ();
 FILLCELL_X1 FILLER_143_818 ();
 FILLCELL_X1 FILLER_143_823 ();
 FILLCELL_X2 FILLER_143_849 ();
 FILLCELL_X4 FILLER_143_855 ();
 FILLCELL_X1 FILLER_143_883 ();
 FILLCELL_X4 FILLER_143_892 ();
 FILLCELL_X4 FILLER_143_918 ();
 FILLCELL_X2 FILLER_143_926 ();
 FILLCELL_X1 FILLER_143_932 ();
 FILLCELL_X2 FILLER_143_936 ();
 FILLCELL_X2 FILLER_143_948 ();
 FILLCELL_X1 FILLER_143_957 ();
 FILLCELL_X1 FILLER_143_971 ();
 FILLCELL_X2 FILLER_143_989 ();
 FILLCELL_X4 FILLER_143_1015 ();
 FILLCELL_X4 FILLER_143_1053 ();
 FILLCELL_X2 FILLER_143_1057 ();
 FILLCELL_X2 FILLER_143_1098 ();
 FILLCELL_X1 FILLER_143_1100 ();
 FILLCELL_X8 FILLER_143_1104 ();
 FILLCELL_X1 FILLER_143_1112 ();
 FILLCELL_X1 FILLER_143_1127 ();
 FILLCELL_X8 FILLER_143_1130 ();
 FILLCELL_X2 FILLER_143_1138 ();
 FILLCELL_X1 FILLER_143_1140 ();
 FILLCELL_X1 FILLER_143_1157 ();
 FILLCELL_X32 FILLER_143_1189 ();
 FILLCELL_X32 FILLER_143_1221 ();
 FILLCELL_X2 FILLER_143_1253 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X8 FILLER_144_65 ();
 FILLCELL_X4 FILLER_144_73 ();
 FILLCELL_X2 FILLER_144_77 ();
 FILLCELL_X4 FILLER_144_84 ();
 FILLCELL_X1 FILLER_144_88 ();
 FILLCELL_X4 FILLER_144_109 ();
 FILLCELL_X1 FILLER_144_113 ();
 FILLCELL_X8 FILLER_144_142 ();
 FILLCELL_X1 FILLER_144_150 ();
 FILLCELL_X4 FILLER_144_158 ();
 FILLCELL_X2 FILLER_144_162 ();
 FILLCELL_X4 FILLER_144_178 ();
 FILLCELL_X2 FILLER_144_182 ();
 FILLCELL_X16 FILLER_144_191 ();
 FILLCELL_X8 FILLER_144_207 ();
 FILLCELL_X4 FILLER_144_215 ();
 FILLCELL_X2 FILLER_144_219 ();
 FILLCELL_X1 FILLER_144_221 ();
 FILLCELL_X1 FILLER_144_229 ();
 FILLCELL_X8 FILLER_144_237 ();
 FILLCELL_X4 FILLER_144_245 ();
 FILLCELL_X2 FILLER_144_249 ();
 FILLCELL_X1 FILLER_144_251 ();
 FILLCELL_X2 FILLER_144_266 ();
 FILLCELL_X1 FILLER_144_268 ();
 FILLCELL_X4 FILLER_144_276 ();
 FILLCELL_X1 FILLER_144_280 ();
 FILLCELL_X2 FILLER_144_288 ();
 FILLCELL_X4 FILLER_144_311 ();
 FILLCELL_X8 FILLER_144_340 ();
 FILLCELL_X2 FILLER_144_348 ();
 FILLCELL_X8 FILLER_144_357 ();
 FILLCELL_X1 FILLER_144_365 ();
 FILLCELL_X4 FILLER_144_374 ();
 FILLCELL_X2 FILLER_144_378 ();
 FILLCELL_X8 FILLER_144_384 ();
 FILLCELL_X1 FILLER_144_392 ();
 FILLCELL_X4 FILLER_144_401 ();
 FILLCELL_X2 FILLER_144_405 ();
 FILLCELL_X4 FILLER_144_441 ();
 FILLCELL_X1 FILLER_144_445 ();
 FILLCELL_X2 FILLER_144_476 ();
 FILLCELL_X1 FILLER_144_478 ();
 FILLCELL_X4 FILLER_144_486 ();
 FILLCELL_X2 FILLER_144_490 ();
 FILLCELL_X1 FILLER_144_492 ();
 FILLCELL_X8 FILLER_144_500 ();
 FILLCELL_X1 FILLER_144_508 ();
 FILLCELL_X1 FILLER_144_517 ();
 FILLCELL_X8 FILLER_144_545 ();
 FILLCELL_X1 FILLER_144_553 ();
 FILLCELL_X32 FILLER_144_581 ();
 FILLCELL_X16 FILLER_144_613 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X4 FILLER_144_696 ();
 FILLCELL_X16 FILLER_144_716 ();
 FILLCELL_X8 FILLER_144_736 ();
 FILLCELL_X4 FILLER_144_744 ();
 FILLCELL_X1 FILLER_144_748 ();
 FILLCELL_X16 FILLER_144_753 ();
 FILLCELL_X1 FILLER_144_771 ();
 FILLCELL_X8 FILLER_144_790 ();
 FILLCELL_X2 FILLER_144_798 ();
 FILLCELL_X1 FILLER_144_800 ();
 FILLCELL_X4 FILLER_144_811 ();
 FILLCELL_X2 FILLER_144_815 ();
 FILLCELL_X1 FILLER_144_827 ();
 FILLCELL_X1 FILLER_144_877 ();
 FILLCELL_X2 FILLER_144_911 ();
 FILLCELL_X4 FILLER_144_925 ();
 FILLCELL_X1 FILLER_144_929 ();
 FILLCELL_X2 FILLER_144_961 ();
 FILLCELL_X4 FILLER_144_973 ();
 FILLCELL_X1 FILLER_144_977 ();
 FILLCELL_X4 FILLER_144_1023 ();
 FILLCELL_X1 FILLER_144_1027 ();
 FILLCELL_X4 FILLER_144_1076 ();
 FILLCELL_X2 FILLER_144_1080 ();
 FILLCELL_X4 FILLER_144_1085 ();
 FILLCELL_X2 FILLER_144_1089 ();
 FILLCELL_X1 FILLER_144_1091 ();
 FILLCELL_X1 FILLER_144_1126 ();
 FILLCELL_X2 FILLER_144_1129 ();
 FILLCELL_X1 FILLER_144_1131 ();
 FILLCELL_X8 FILLER_144_1144 ();
 FILLCELL_X2 FILLER_144_1152 ();
 FILLCELL_X32 FILLER_144_1187 ();
 FILLCELL_X32 FILLER_144_1219 ();
 FILLCELL_X4 FILLER_144_1251 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X8 FILLER_145_65 ();
 FILLCELL_X4 FILLER_145_73 ();
 FILLCELL_X1 FILLER_145_77 ();
 FILLCELL_X4 FILLER_145_98 ();
 FILLCELL_X1 FILLER_145_102 ();
 FILLCELL_X8 FILLER_145_137 ();
 FILLCELL_X4 FILLER_145_152 ();
 FILLCELL_X2 FILLER_145_156 ();
 FILLCELL_X1 FILLER_145_158 ();
 FILLCELL_X4 FILLER_145_179 ();
 FILLCELL_X2 FILLER_145_183 ();
 FILLCELL_X4 FILLER_145_192 ();
 FILLCELL_X2 FILLER_145_196 ();
 FILLCELL_X1 FILLER_145_198 ();
 FILLCELL_X2 FILLER_145_240 ();
 FILLCELL_X8 FILLER_145_249 ();
 FILLCELL_X4 FILLER_145_264 ();
 FILLCELL_X8 FILLER_145_302 ();
 FILLCELL_X1 FILLER_145_330 ();
 FILLCELL_X1 FILLER_145_338 ();
 FILLCELL_X1 FILLER_145_346 ();
 FILLCELL_X4 FILLER_145_367 ();
 FILLCELL_X2 FILLER_145_371 ();
 FILLCELL_X2 FILLER_145_400 ();
 FILLCELL_X8 FILLER_145_412 ();
 FILLCELL_X4 FILLER_145_420 ();
 FILLCELL_X1 FILLER_145_424 ();
 FILLCELL_X32 FILLER_145_432 ();
 FILLCELL_X2 FILLER_145_464 ();
 FILLCELL_X8 FILLER_145_469 ();
 FILLCELL_X1 FILLER_145_477 ();
 FILLCELL_X2 FILLER_145_519 ();
 FILLCELL_X1 FILLER_145_521 ();
 FILLCELL_X2 FILLER_145_529 ();
 FILLCELL_X2 FILLER_145_545 ();
 FILLCELL_X1 FILLER_145_547 ();
 FILLCELL_X2 FILLER_145_574 ();
 FILLCELL_X32 FILLER_145_583 ();
 FILLCELL_X32 FILLER_145_615 ();
 FILLCELL_X32 FILLER_145_647 ();
 FILLCELL_X16 FILLER_145_679 ();
 FILLCELL_X4 FILLER_145_695 ();
 FILLCELL_X2 FILLER_145_699 ();
 FILLCELL_X1 FILLER_145_701 ();
 FILLCELL_X1 FILLER_145_708 ();
 FILLCELL_X2 FILLER_145_715 ();
 FILLCELL_X2 FILLER_145_721 ();
 FILLCELL_X1 FILLER_145_739 ();
 FILLCELL_X4 FILLER_145_756 ();
 FILLCELL_X2 FILLER_145_760 ();
 FILLCELL_X4 FILLER_145_778 ();
 FILLCELL_X2 FILLER_145_782 ();
 FILLCELL_X1 FILLER_145_784 ();
 FILLCELL_X4 FILLER_145_814 ();
 FILLCELL_X4 FILLER_145_847 ();
 FILLCELL_X1 FILLER_145_851 ();
 FILLCELL_X1 FILLER_145_857 ();
 FILLCELL_X1 FILLER_145_873 ();
 FILLCELL_X2 FILLER_145_880 ();
 FILLCELL_X1 FILLER_145_882 ();
 FILLCELL_X4 FILLER_145_919 ();
 FILLCELL_X1 FILLER_145_937 ();
 FILLCELL_X2 FILLER_145_955 ();
 FILLCELL_X1 FILLER_145_957 ();
 FILLCELL_X4 FILLER_145_961 ();
 FILLCELL_X1 FILLER_145_965 ();
 FILLCELL_X2 FILLER_145_968 ();
 FILLCELL_X8 FILLER_145_972 ();
 FILLCELL_X4 FILLER_145_980 ();
 FILLCELL_X8 FILLER_145_1017 ();
 FILLCELL_X4 FILLER_145_1025 ();
 FILLCELL_X1 FILLER_145_1029 ();
 FILLCELL_X1 FILLER_145_1043 ();
 FILLCELL_X4 FILLER_145_1047 ();
 FILLCELL_X1 FILLER_145_1051 ();
 FILLCELL_X4 FILLER_145_1057 ();
 FILLCELL_X2 FILLER_145_1061 ();
 FILLCELL_X4 FILLER_145_1068 ();
 FILLCELL_X2 FILLER_145_1072 ();
 FILLCELL_X2 FILLER_145_1076 ();
 FILLCELL_X2 FILLER_145_1081 ();
 FILLCELL_X4 FILLER_145_1093 ();
 FILLCELL_X1 FILLER_145_1097 ();
 FILLCELL_X32 FILLER_145_1199 ();
 FILLCELL_X16 FILLER_145_1231 ();
 FILLCELL_X2 FILLER_145_1247 ();
 FILLCELL_X1 FILLER_145_1251 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X16 FILLER_146_65 ();
 FILLCELL_X8 FILLER_146_81 ();
 FILLCELL_X2 FILLER_146_89 ();
 FILLCELL_X1 FILLER_146_91 ();
 FILLCELL_X4 FILLER_146_99 ();
 FILLCELL_X2 FILLER_146_103 ();
 FILLCELL_X1 FILLER_146_105 ();
 FILLCELL_X4 FILLER_146_117 ();
 FILLCELL_X2 FILLER_146_128 ();
 FILLCELL_X1 FILLER_146_130 ();
 FILLCELL_X1 FILLER_146_138 ();
 FILLCELL_X2 FILLER_146_146 ();
 FILLCELL_X1 FILLER_146_148 ();
 FILLCELL_X8 FILLER_146_156 ();
 FILLCELL_X4 FILLER_146_164 ();
 FILLCELL_X2 FILLER_146_168 ();
 FILLCELL_X1 FILLER_146_170 ();
 FILLCELL_X4 FILLER_146_178 ();
 FILLCELL_X2 FILLER_146_182 ();
 FILLCELL_X1 FILLER_146_184 ();
 FILLCELL_X4 FILLER_146_206 ();
 FILLCELL_X2 FILLER_146_210 ();
 FILLCELL_X1 FILLER_146_259 ();
 FILLCELL_X1 FILLER_146_267 ();
 FILLCELL_X1 FILLER_146_275 ();
 FILLCELL_X2 FILLER_146_296 ();
 FILLCELL_X1 FILLER_146_298 ();
 FILLCELL_X8 FILLER_146_306 ();
 FILLCELL_X8 FILLER_146_321 ();
 FILLCELL_X2 FILLER_146_329 ();
 FILLCELL_X1 FILLER_146_331 ();
 FILLCELL_X4 FILLER_146_339 ();
 FILLCELL_X1 FILLER_146_343 ();
 FILLCELL_X2 FILLER_146_351 ();
 FILLCELL_X2 FILLER_146_360 ();
 FILLCELL_X4 FILLER_146_389 ();
 FILLCELL_X1 FILLER_146_393 ();
 FILLCELL_X2 FILLER_146_408 ();
 FILLCELL_X8 FILLER_146_413 ();
 FILLCELL_X1 FILLER_146_421 ();
 FILLCELL_X2 FILLER_146_456 ();
 FILLCELL_X4 FILLER_146_472 ();
 FILLCELL_X2 FILLER_146_476 ();
 FILLCELL_X1 FILLER_146_478 ();
 FILLCELL_X1 FILLER_146_497 ();
 FILLCELL_X4 FILLER_146_502 ();
 FILLCELL_X2 FILLER_146_506 ();
 FILLCELL_X1 FILLER_146_508 ();
 FILLCELL_X4 FILLER_146_536 ();
 FILLCELL_X1 FILLER_146_547 ();
 FILLCELL_X2 FILLER_146_555 ();
 FILLCELL_X4 FILLER_146_564 ();
 FILLCELL_X2 FILLER_146_568 ();
 FILLCELL_X32 FILLER_146_590 ();
 FILLCELL_X8 FILLER_146_622 ();
 FILLCELL_X1 FILLER_146_630 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X2 FILLER_146_696 ();
 FILLCELL_X4 FILLER_146_724 ();
 FILLCELL_X1 FILLER_146_728 ();
 FILLCELL_X2 FILLER_146_743 ();
 FILLCELL_X8 FILLER_146_761 ();
 FILLCELL_X4 FILLER_146_769 ();
 FILLCELL_X2 FILLER_146_773 ();
 FILLCELL_X1 FILLER_146_775 ();
 FILLCELL_X8 FILLER_146_778 ();
 FILLCELL_X1 FILLER_146_786 ();
 FILLCELL_X2 FILLER_146_799 ();
 FILLCELL_X1 FILLER_146_805 ();
 FILLCELL_X1 FILLER_146_818 ();
 FILLCELL_X4 FILLER_146_825 ();
 FILLCELL_X2 FILLER_146_829 ();
 FILLCELL_X1 FILLER_146_831 ();
 FILLCELL_X4 FILLER_146_838 ();
 FILLCELL_X1 FILLER_146_842 ();
 FILLCELL_X1 FILLER_146_868 ();
 FILLCELL_X4 FILLER_146_876 ();
 FILLCELL_X2 FILLER_146_884 ();
 FILLCELL_X1 FILLER_146_901 ();
 FILLCELL_X8 FILLER_146_907 ();
 FILLCELL_X2 FILLER_146_915 ();
 FILLCELL_X1 FILLER_146_917 ();
 FILLCELL_X1 FILLER_146_939 ();
 FILLCELL_X1 FILLER_146_944 ();
 FILLCELL_X8 FILLER_146_993 ();
 FILLCELL_X4 FILLER_146_1001 ();
 FILLCELL_X1 FILLER_146_1015 ();
 FILLCELL_X2 FILLER_146_1033 ();
 FILLCELL_X4 FILLER_146_1053 ();
 FILLCELL_X1 FILLER_146_1089 ();
 FILLCELL_X4 FILLER_146_1112 ();
 FILLCELL_X2 FILLER_146_1116 ();
 FILLCELL_X8 FILLER_146_1120 ();
 FILLCELL_X1 FILLER_146_1128 ();
 FILLCELL_X4 FILLER_146_1131 ();
 FILLCELL_X2 FILLER_146_1135 ();
 FILLCELL_X1 FILLER_146_1137 ();
 FILLCELL_X8 FILLER_146_1140 ();
 FILLCELL_X4 FILLER_146_1148 ();
 FILLCELL_X1 FILLER_146_1152 ();
 FILLCELL_X1 FILLER_146_1155 ();
 FILLCELL_X8 FILLER_146_1158 ();
 FILLCELL_X1 FILLER_146_1166 ();
 FILLCELL_X2 FILLER_146_1186 ();
 FILLCELL_X32 FILLER_146_1197 ();
 FILLCELL_X8 FILLER_146_1229 ();
 FILLCELL_X4 FILLER_146_1247 ();
 FILLCELL_X1 FILLER_146_1254 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X8 FILLER_147_65 ();
 FILLCELL_X2 FILLER_147_73 ();
 FILLCELL_X8 FILLER_147_102 ();
 FILLCELL_X4 FILLER_147_110 ();
 FILLCELL_X1 FILLER_147_114 ();
 FILLCELL_X4 FILLER_147_157 ();
 FILLCELL_X2 FILLER_147_181 ();
 FILLCELL_X1 FILLER_147_190 ();
 FILLCELL_X2 FILLER_147_198 ();
 FILLCELL_X1 FILLER_147_200 ();
 FILLCELL_X4 FILLER_147_213 ();
 FILLCELL_X1 FILLER_147_217 ();
 FILLCELL_X2 FILLER_147_225 ();
 FILLCELL_X8 FILLER_147_234 ();
 FILLCELL_X1 FILLER_147_242 ();
 FILLCELL_X16 FILLER_147_264 ();
 FILLCELL_X4 FILLER_147_280 ();
 FILLCELL_X16 FILLER_147_296 ();
 FILLCELL_X4 FILLER_147_312 ();
 FILLCELL_X2 FILLER_147_316 ();
 FILLCELL_X4 FILLER_147_338 ();
 FILLCELL_X2 FILLER_147_342 ();
 FILLCELL_X1 FILLER_147_364 ();
 FILLCELL_X8 FILLER_147_399 ();
 FILLCELL_X4 FILLER_147_407 ();
 FILLCELL_X2 FILLER_147_411 ();
 FILLCELL_X1 FILLER_147_413 ();
 FILLCELL_X1 FILLER_147_427 ();
 FILLCELL_X1 FILLER_147_435 ();
 FILLCELL_X16 FILLER_147_463 ();
 FILLCELL_X2 FILLER_147_479 ();
 FILLCELL_X1 FILLER_147_481 ();
 FILLCELL_X8 FILLER_147_499 ();
 FILLCELL_X2 FILLER_147_507 ();
 FILLCELL_X1 FILLER_147_509 ();
 FILLCELL_X1 FILLER_147_517 ();
 FILLCELL_X2 FILLER_147_546 ();
 FILLCELL_X32 FILLER_147_575 ();
 FILLCELL_X32 FILLER_147_607 ();
 FILLCELL_X32 FILLER_147_639 ();
 FILLCELL_X32 FILLER_147_671 ();
 FILLCELL_X4 FILLER_147_719 ();
 FILLCELL_X1 FILLER_147_723 ();
 FILLCELL_X4 FILLER_147_742 ();
 FILLCELL_X2 FILLER_147_746 ();
 FILLCELL_X4 FILLER_147_750 ();
 FILLCELL_X4 FILLER_147_764 ();
 FILLCELL_X2 FILLER_147_768 ();
 FILLCELL_X1 FILLER_147_770 ();
 FILLCELL_X2 FILLER_147_781 ();
 FILLCELL_X2 FILLER_147_795 ();
 FILLCELL_X4 FILLER_147_815 ();
 FILLCELL_X4 FILLER_147_855 ();
 FILLCELL_X1 FILLER_147_859 ();
 FILLCELL_X1 FILLER_147_924 ();
 FILLCELL_X1 FILLER_147_975 ();
 FILLCELL_X2 FILLER_147_980 ();
 FILLCELL_X1 FILLER_147_982 ();
 FILLCELL_X1 FILLER_147_992 ();
 FILLCELL_X1 FILLER_147_1009 ();
 FILLCELL_X8 FILLER_147_1012 ();
 FILLCELL_X4 FILLER_147_1020 ();
 FILLCELL_X1 FILLER_147_1024 ();
 FILLCELL_X16 FILLER_147_1028 ();
 FILLCELL_X16 FILLER_147_1059 ();
 FILLCELL_X4 FILLER_147_1075 ();
 FILLCELL_X1 FILLER_147_1079 ();
 FILLCELL_X16 FILLER_147_1086 ();
 FILLCELL_X2 FILLER_147_1102 ();
 FILLCELL_X1 FILLER_147_1130 ();
 FILLCELL_X16 FILLER_147_1157 ();
 FILLCELL_X4 FILLER_147_1173 ();
 FILLCELL_X2 FILLER_147_1177 ();
 FILLCELL_X1 FILLER_147_1179 ();
 FILLCELL_X32 FILLER_147_1201 ();
 FILLCELL_X8 FILLER_147_1233 ();
 FILLCELL_X2 FILLER_147_1241 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X1 FILLER_148_124 ();
 FILLCELL_X1 FILLER_148_159 ();
 FILLCELL_X2 FILLER_148_206 ();
 FILLCELL_X2 FILLER_148_215 ();
 FILLCELL_X2 FILLER_148_265 ();
 FILLCELL_X2 FILLER_148_287 ();
 FILLCELL_X1 FILLER_148_289 ();
 FILLCELL_X4 FILLER_148_311 ();
 FILLCELL_X8 FILLER_148_336 ();
 FILLCELL_X4 FILLER_148_344 ();
 FILLCELL_X2 FILLER_148_348 ();
 FILLCELL_X1 FILLER_148_350 ();
 FILLCELL_X4 FILLER_148_358 ();
 FILLCELL_X4 FILLER_148_369 ();
 FILLCELL_X2 FILLER_148_394 ();
 FILLCELL_X2 FILLER_148_399 ();
 FILLCELL_X8 FILLER_148_440 ();
 FILLCELL_X4 FILLER_148_448 ();
 FILLCELL_X2 FILLER_148_479 ();
 FILLCELL_X1 FILLER_148_481 ();
 FILLCELL_X2 FILLER_148_509 ();
 FILLCELL_X4 FILLER_148_531 ();
 FILLCELL_X4 FILLER_148_542 ();
 FILLCELL_X2 FILLER_148_553 ();
 FILLCELL_X1 FILLER_148_555 ();
 FILLCELL_X32 FILLER_148_583 ();
 FILLCELL_X16 FILLER_148_615 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X8 FILLER_148_696 ();
 FILLCELL_X2 FILLER_148_704 ();
 FILLCELL_X4 FILLER_148_712 ();
 FILLCELL_X2 FILLER_148_716 ();
 FILLCELL_X8 FILLER_148_720 ();
 FILLCELL_X1 FILLER_148_728 ();
 FILLCELL_X4 FILLER_148_767 ();
 FILLCELL_X8 FILLER_148_801 ();
 FILLCELL_X2 FILLER_148_809 ();
 FILLCELL_X4 FILLER_148_813 ();
 FILLCELL_X4 FILLER_148_828 ();
 FILLCELL_X2 FILLER_148_832 ();
 FILLCELL_X2 FILLER_148_836 ();
 FILLCELL_X1 FILLER_148_838 ();
 FILLCELL_X1 FILLER_148_843 ();
 FILLCELL_X8 FILLER_148_864 ();
 FILLCELL_X8 FILLER_148_876 ();
 FILLCELL_X4 FILLER_148_884 ();
 FILLCELL_X8 FILLER_148_892 ();
 FILLCELL_X4 FILLER_148_900 ();
 FILLCELL_X1 FILLER_148_904 ();
 FILLCELL_X8 FILLER_148_909 ();
 FILLCELL_X4 FILLER_148_917 ();
 FILLCELL_X1 FILLER_148_921 ();
 FILLCELL_X8 FILLER_148_928 ();
 FILLCELL_X4 FILLER_148_936 ();
 FILLCELL_X2 FILLER_148_940 ();
 FILLCELL_X8 FILLER_148_946 ();
 FILLCELL_X2 FILLER_148_954 ();
 FILLCELL_X1 FILLER_148_956 ();
 FILLCELL_X1 FILLER_148_959 ();
 FILLCELL_X1 FILLER_148_969 ();
 FILLCELL_X8 FILLER_148_1002 ();
 FILLCELL_X1 FILLER_148_1010 ();
 FILLCELL_X4 FILLER_148_1035 ();
 FILLCELL_X2 FILLER_148_1039 ();
 FILLCELL_X4 FILLER_148_1073 ();
 FILLCELL_X8 FILLER_148_1085 ();
 FILLCELL_X16 FILLER_148_1099 ();
 FILLCELL_X4 FILLER_148_1115 ();
 FILLCELL_X1 FILLER_148_1119 ();
 FILLCELL_X1 FILLER_148_1122 ();
 FILLCELL_X1 FILLER_148_1125 ();
 FILLCELL_X1 FILLER_148_1179 ();
 FILLCELL_X32 FILLER_148_1200 ();
 FILLCELL_X16 FILLER_148_1232 ();
 FILLCELL_X4 FILLER_148_1248 ();
 FILLCELL_X2 FILLER_148_1252 ();
 FILLCELL_X1 FILLER_148_1254 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X16 FILLER_149_97 ();
 FILLCELL_X4 FILLER_149_113 ();
 FILLCELL_X2 FILLER_149_149 ();
 FILLCELL_X8 FILLER_149_174 ();
 FILLCELL_X2 FILLER_149_182 ();
 FILLCELL_X1 FILLER_149_184 ();
 FILLCELL_X1 FILLER_149_206 ();
 FILLCELL_X4 FILLER_149_262 ();
 FILLCELL_X2 FILLER_149_266 ();
 FILLCELL_X4 FILLER_149_275 ();
 FILLCELL_X1 FILLER_149_279 ();
 FILLCELL_X1 FILLER_149_294 ();
 FILLCELL_X8 FILLER_149_335 ();
 FILLCELL_X1 FILLER_149_363 ();
 FILLCELL_X16 FILLER_149_378 ();
 FILLCELL_X2 FILLER_149_394 ();
 FILLCELL_X16 FILLER_149_399 ();
 FILLCELL_X1 FILLER_149_435 ();
 FILLCELL_X1 FILLER_149_445 ();
 FILLCELL_X4 FILLER_149_453 ();
 FILLCELL_X2 FILLER_149_457 ();
 FILLCELL_X4 FILLER_149_464 ();
 FILLCELL_X2 FILLER_149_468 ();
 FILLCELL_X1 FILLER_149_470 ();
 FILLCELL_X4 FILLER_149_478 ();
 FILLCELL_X8 FILLER_149_489 ();
 FILLCELL_X1 FILLER_149_504 ();
 FILLCELL_X4 FILLER_149_532 ();
 FILLCELL_X2 FILLER_149_536 ();
 FILLCELL_X1 FILLER_149_538 ();
 FILLCELL_X32 FILLER_149_559 ();
 FILLCELL_X32 FILLER_149_591 ();
 FILLCELL_X32 FILLER_149_623 ();
 FILLCELL_X32 FILLER_149_655 ();
 FILLCELL_X16 FILLER_149_687 ();
 FILLCELL_X2 FILLER_149_709 ();
 FILLCELL_X4 FILLER_149_743 ();
 FILLCELL_X4 FILLER_149_765 ();
 FILLCELL_X2 FILLER_149_769 ();
 FILLCELL_X1 FILLER_149_771 ();
 FILLCELL_X1 FILLER_149_774 ();
 FILLCELL_X4 FILLER_149_821 ();
 FILLCELL_X2 FILLER_149_863 ();
 FILLCELL_X1 FILLER_149_865 ();
 FILLCELL_X4 FILLER_149_932 ();
 FILLCELL_X1 FILLER_149_936 ();
 FILLCELL_X1 FILLER_149_953 ();
 FILLCELL_X8 FILLER_149_982 ();
 FILLCELL_X2 FILLER_149_990 ();
 FILLCELL_X1 FILLER_149_992 ();
 FILLCELL_X2 FILLER_149_1030 ();
 FILLCELL_X2 FILLER_149_1035 ();
 FILLCELL_X8 FILLER_149_1053 ();
 FILLCELL_X1 FILLER_149_1120 ();
 FILLCELL_X16 FILLER_149_1138 ();
 FILLCELL_X4 FILLER_149_1154 ();
 FILLCELL_X2 FILLER_149_1158 ();
 FILLCELL_X1 FILLER_149_1160 ();
 FILLCELL_X1 FILLER_149_1163 ();
 FILLCELL_X32 FILLER_149_1203 ();
 FILLCELL_X16 FILLER_149_1235 ();
 FILLCELL_X4 FILLER_149_1251 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X4 FILLER_150_97 ();
 FILLCELL_X2 FILLER_150_101 ();
 FILLCELL_X32 FILLER_150_130 ();
 FILLCELL_X16 FILLER_150_162 ();
 FILLCELL_X1 FILLER_150_178 ();
 FILLCELL_X8 FILLER_150_206 ();
 FILLCELL_X4 FILLER_150_214 ();
 FILLCELL_X2 FILLER_150_218 ();
 FILLCELL_X16 FILLER_150_227 ();
 FILLCELL_X8 FILLER_150_243 ();
 FILLCELL_X4 FILLER_150_251 ();
 FILLCELL_X1 FILLER_150_255 ();
 FILLCELL_X1 FILLER_150_303 ();
 FILLCELL_X4 FILLER_150_331 ();
 FILLCELL_X2 FILLER_150_335 ();
 FILLCELL_X2 FILLER_150_342 ();
 FILLCELL_X8 FILLER_150_351 ();
 FILLCELL_X1 FILLER_150_359 ();
 FILLCELL_X4 FILLER_150_374 ();
 FILLCELL_X2 FILLER_150_378 ();
 FILLCELL_X1 FILLER_150_380 ();
 FILLCELL_X4 FILLER_150_388 ();
 FILLCELL_X1 FILLER_150_392 ();
 FILLCELL_X4 FILLER_150_414 ();
 FILLCELL_X2 FILLER_150_418 ();
 FILLCELL_X1 FILLER_150_420 ();
 FILLCELL_X1 FILLER_150_428 ();
 FILLCELL_X2 FILLER_150_436 ();
 FILLCELL_X2 FILLER_150_445 ();
 FILLCELL_X1 FILLER_150_447 ();
 FILLCELL_X1 FILLER_150_455 ();
 FILLCELL_X2 FILLER_150_476 ();
 FILLCELL_X1 FILLER_150_478 ();
 FILLCELL_X8 FILLER_150_486 ();
 FILLCELL_X4 FILLER_150_494 ();
 FILLCELL_X32 FILLER_150_525 ();
 FILLCELL_X32 FILLER_150_557 ();
 FILLCELL_X32 FILLER_150_589 ();
 FILLCELL_X8 FILLER_150_621 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X8 FILLER_150_696 ();
 FILLCELL_X1 FILLER_150_710 ();
 FILLCELL_X4 FILLER_150_717 ();
 FILLCELL_X1 FILLER_150_721 ();
 FILLCELL_X16 FILLER_150_734 ();
 FILLCELL_X8 FILLER_150_750 ();
 FILLCELL_X2 FILLER_150_758 ();
 FILLCELL_X1 FILLER_150_760 ();
 FILLCELL_X2 FILLER_150_779 ();
 FILLCELL_X1 FILLER_150_781 ();
 FILLCELL_X4 FILLER_150_784 ();
 FILLCELL_X2 FILLER_150_788 ();
 FILLCELL_X4 FILLER_150_792 ();
 FILLCELL_X2 FILLER_150_796 ();
 FILLCELL_X16 FILLER_150_800 ();
 FILLCELL_X8 FILLER_150_816 ();
 FILLCELL_X1 FILLER_150_824 ();
 FILLCELL_X8 FILLER_150_827 ();
 FILLCELL_X1 FILLER_150_835 ();
 FILLCELL_X4 FILLER_150_846 ();
 FILLCELL_X2 FILLER_150_850 ();
 FILLCELL_X2 FILLER_150_854 ();
 FILLCELL_X16 FILLER_150_858 ();
 FILLCELL_X4 FILLER_150_874 ();
 FILLCELL_X1 FILLER_150_882 ();
 FILLCELL_X4 FILLER_150_886 ();
 FILLCELL_X2 FILLER_150_890 ();
 FILLCELL_X8 FILLER_150_896 ();
 FILLCELL_X1 FILLER_150_904 ();
 FILLCELL_X8 FILLER_150_907 ();
 FILLCELL_X2 FILLER_150_915 ();
 FILLCELL_X2 FILLER_150_919 ();
 FILLCELL_X1 FILLER_150_921 ();
 FILLCELL_X4 FILLER_150_942 ();
 FILLCELL_X1 FILLER_150_946 ();
 FILLCELL_X4 FILLER_150_949 ();
 FILLCELL_X1 FILLER_150_974 ();
 FILLCELL_X4 FILLER_150_1007 ();
 FILLCELL_X1 FILLER_150_1011 ();
 FILLCELL_X4 FILLER_150_1015 ();
 FILLCELL_X8 FILLER_150_1041 ();
 FILLCELL_X1 FILLER_150_1049 ();
 FILLCELL_X4 FILLER_150_1073 ();
 FILLCELL_X2 FILLER_150_1077 ();
 FILLCELL_X1 FILLER_150_1079 ();
 FILLCELL_X4 FILLER_150_1091 ();
 FILLCELL_X1 FILLER_150_1095 ();
 FILLCELL_X1 FILLER_150_1099 ();
 FILLCELL_X1 FILLER_150_1108 ();
 FILLCELL_X1 FILLER_150_1111 ();
 FILLCELL_X4 FILLER_150_1115 ();
 FILLCELL_X16 FILLER_150_1147 ();
 FILLCELL_X4 FILLER_150_1173 ();
 FILLCELL_X32 FILLER_150_1203 ();
 FILLCELL_X16 FILLER_150_1235 ();
 FILLCELL_X4 FILLER_150_1251 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X4 FILLER_151_97 ();
 FILLCELL_X2 FILLER_151_101 ();
 FILLCELL_X1 FILLER_151_103 ();
 FILLCELL_X2 FILLER_151_131 ();
 FILLCELL_X8 FILLER_151_160 ();
 FILLCELL_X16 FILLER_151_195 ();
 FILLCELL_X8 FILLER_151_211 ();
 FILLCELL_X2 FILLER_151_219 ();
 FILLCELL_X16 FILLER_151_248 ();
 FILLCELL_X4 FILLER_151_271 ();
 FILLCELL_X1 FILLER_151_275 ();
 FILLCELL_X32 FILLER_151_296 ();
 FILLCELL_X2 FILLER_151_328 ();
 FILLCELL_X1 FILLER_151_330 ();
 FILLCELL_X4 FILLER_151_375 ();
 FILLCELL_X1 FILLER_151_399 ();
 FILLCELL_X2 FILLER_151_414 ();
 FILLCELL_X1 FILLER_151_416 ();
 FILLCELL_X16 FILLER_151_451 ();
 FILLCELL_X4 FILLER_151_467 ();
 FILLCELL_X4 FILLER_151_492 ();
 FILLCELL_X2 FILLER_151_496 ();
 FILLCELL_X32 FILLER_151_530 ();
 FILLCELL_X32 FILLER_151_562 ();
 FILLCELL_X32 FILLER_151_594 ();
 FILLCELL_X32 FILLER_151_626 ();
 FILLCELL_X32 FILLER_151_658 ();
 FILLCELL_X8 FILLER_151_690 ();
 FILLCELL_X4 FILLER_151_698 ();
 FILLCELL_X2 FILLER_151_702 ();
 FILLCELL_X1 FILLER_151_704 ();
 FILLCELL_X1 FILLER_151_711 ();
 FILLCELL_X1 FILLER_151_718 ();
 FILLCELL_X8 FILLER_151_725 ();
 FILLCELL_X2 FILLER_151_749 ();
 FILLCELL_X2 FILLER_151_767 ();
 FILLCELL_X1 FILLER_151_769 ();
 FILLCELL_X8 FILLER_151_773 ();
 FILLCELL_X2 FILLER_151_781 ();
 FILLCELL_X2 FILLER_151_825 ();
 FILLCELL_X1 FILLER_151_845 ();
 FILLCELL_X2 FILLER_151_848 ();
 FILLCELL_X4 FILLER_151_860 ();
 FILLCELL_X2 FILLER_151_886 ();
 FILLCELL_X1 FILLER_151_888 ();
 FILLCELL_X1 FILLER_151_899 ();
 FILLCELL_X8 FILLER_151_913 ();
 FILLCELL_X1 FILLER_151_921 ();
 FILLCELL_X1 FILLER_151_924 ();
 FILLCELL_X2 FILLER_151_929 ();
 FILLCELL_X4 FILLER_151_933 ();
 FILLCELL_X1 FILLER_151_937 ();
 FILLCELL_X8 FILLER_151_948 ();
 FILLCELL_X1 FILLER_151_956 ();
 FILLCELL_X8 FILLER_151_960 ();
 FILLCELL_X2 FILLER_151_968 ();
 FILLCELL_X1 FILLER_151_970 ();
 FILLCELL_X2 FILLER_151_975 ();
 FILLCELL_X8 FILLER_151_980 ();
 FILLCELL_X2 FILLER_151_990 ();
 FILLCELL_X1 FILLER_151_1010 ();
 FILLCELL_X8 FILLER_151_1013 ();
 FILLCELL_X2 FILLER_151_1021 ();
 FILLCELL_X1 FILLER_151_1026 ();
 FILLCELL_X2 FILLER_151_1030 ();
 FILLCELL_X2 FILLER_151_1048 ();
 FILLCELL_X4 FILLER_151_1062 ();
 FILLCELL_X4 FILLER_151_1068 ();
 FILLCELL_X2 FILLER_151_1072 ();
 FILLCELL_X1 FILLER_151_1076 ();
 FILLCELL_X4 FILLER_151_1113 ();
 FILLCELL_X1 FILLER_151_1117 ();
 FILLCELL_X2 FILLER_151_1120 ();
 FILLCELL_X1 FILLER_151_1132 ();
 FILLCELL_X1 FILLER_151_1135 ();
 FILLCELL_X1 FILLER_151_1146 ();
 FILLCELL_X2 FILLER_151_1150 ();
 FILLCELL_X8 FILLER_151_1157 ();
 FILLCELL_X4 FILLER_151_1165 ();
 FILLCELL_X32 FILLER_151_1190 ();
 FILLCELL_X32 FILLER_151_1222 ();
 FILLCELL_X1 FILLER_151_1254 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X16 FILLER_152_97 ();
 FILLCELL_X8 FILLER_152_113 ();
 FILLCELL_X32 FILLER_152_148 ();
 FILLCELL_X8 FILLER_152_180 ();
 FILLCELL_X2 FILLER_152_188 ();
 FILLCELL_X1 FILLER_152_190 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X16 FILLER_152_257 ();
 FILLCELL_X4 FILLER_152_273 ();
 FILLCELL_X1 FILLER_152_277 ();
 FILLCELL_X4 FILLER_152_285 ();
 FILLCELL_X2 FILLER_152_289 ();
 FILLCELL_X8 FILLER_152_318 ();
 FILLCELL_X4 FILLER_152_326 ();
 FILLCELL_X2 FILLER_152_330 ();
 FILLCELL_X1 FILLER_152_332 ();
 FILLCELL_X2 FILLER_152_360 ();
 FILLCELL_X1 FILLER_152_362 ();
 FILLCELL_X4 FILLER_152_370 ();
 FILLCELL_X1 FILLER_152_374 ();
 FILLCELL_X4 FILLER_152_403 ();
 FILLCELL_X2 FILLER_152_407 ();
 FILLCELL_X1 FILLER_152_409 ();
 FILLCELL_X2 FILLER_152_450 ();
 FILLCELL_X8 FILLER_152_472 ();
 FILLCELL_X4 FILLER_152_480 ();
 FILLCELL_X32 FILLER_152_511 ();
 FILLCELL_X32 FILLER_152_543 ();
 FILLCELL_X32 FILLER_152_575 ();
 FILLCELL_X16 FILLER_152_607 ();
 FILLCELL_X8 FILLER_152_623 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X1 FILLER_152_696 ();
 FILLCELL_X2 FILLER_152_715 ();
 FILLCELL_X8 FILLER_152_721 ();
 FILLCELL_X4 FILLER_152_729 ();
 FILLCELL_X8 FILLER_152_749 ();
 FILLCELL_X4 FILLER_152_757 ();
 FILLCELL_X2 FILLER_152_761 ();
 FILLCELL_X2 FILLER_152_771 ();
 FILLCELL_X1 FILLER_152_794 ();
 FILLCELL_X4 FILLER_152_797 ();
 FILLCELL_X2 FILLER_152_803 ();
 FILLCELL_X1 FILLER_152_805 ();
 FILLCELL_X4 FILLER_152_826 ();
 FILLCELL_X1 FILLER_152_830 ();
 FILLCELL_X8 FILLER_152_833 ();
 FILLCELL_X1 FILLER_152_841 ();
 FILLCELL_X8 FILLER_152_874 ();
 FILLCELL_X1 FILLER_152_920 ();
 FILLCELL_X2 FILLER_152_966 ();
 FILLCELL_X8 FILLER_152_990 ();
 FILLCELL_X2 FILLER_152_998 ();
 FILLCELL_X1 FILLER_152_1000 ();
 FILLCELL_X2 FILLER_152_1003 ();
 FILLCELL_X8 FILLER_152_1037 ();
 FILLCELL_X4 FILLER_152_1045 ();
 FILLCELL_X4 FILLER_152_1097 ();
 FILLCELL_X2 FILLER_152_1101 ();
 FILLCELL_X4 FILLER_152_1119 ();
 FILLCELL_X4 FILLER_152_1135 ();
 FILLCELL_X4 FILLER_152_1171 ();
 FILLCELL_X2 FILLER_152_1175 ();
 FILLCELL_X2 FILLER_152_1181 ();
 FILLCELL_X1 FILLER_152_1183 ();
 FILLCELL_X32 FILLER_152_1191 ();
 FILLCELL_X32 FILLER_152_1223 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X16 FILLER_153_161 ();
 FILLCELL_X2 FILLER_153_177 ();
 FILLCELL_X1 FILLER_153_179 ();
 FILLCELL_X1 FILLER_153_207 ();
 FILLCELL_X32 FILLER_153_228 ();
 FILLCELL_X32 FILLER_153_260 ();
 FILLCELL_X32 FILLER_153_292 ();
 FILLCELL_X16 FILLER_153_324 ();
 FILLCELL_X4 FILLER_153_340 ();
 FILLCELL_X1 FILLER_153_344 ();
 FILLCELL_X1 FILLER_153_372 ();
 FILLCELL_X4 FILLER_153_380 ();
 FILLCELL_X2 FILLER_153_384 ();
 FILLCELL_X4 FILLER_153_413 ();
 FILLCELL_X1 FILLER_153_417 ();
 FILLCELL_X8 FILLER_153_425 ();
 FILLCELL_X2 FILLER_153_433 ();
 FILLCELL_X8 FILLER_153_442 ();
 FILLCELL_X2 FILLER_153_450 ();
 FILLCELL_X4 FILLER_153_459 ();
 FILLCELL_X2 FILLER_153_463 ();
 FILLCELL_X1 FILLER_153_465 ();
 FILLCELL_X32 FILLER_153_493 ();
 FILLCELL_X32 FILLER_153_525 ();
 FILLCELL_X32 FILLER_153_557 ();
 FILLCELL_X32 FILLER_153_589 ();
 FILLCELL_X32 FILLER_153_621 ();
 FILLCELL_X32 FILLER_153_653 ();
 FILLCELL_X16 FILLER_153_685 ();
 FILLCELL_X8 FILLER_153_701 ();
 FILLCELL_X1 FILLER_153_709 ();
 FILLCELL_X4 FILLER_153_726 ();
 FILLCELL_X4 FILLER_153_732 ();
 FILLCELL_X1 FILLER_153_738 ();
 FILLCELL_X2 FILLER_153_741 ();
 FILLCELL_X1 FILLER_153_743 ();
 FILLCELL_X2 FILLER_153_760 ();
 FILLCELL_X1 FILLER_153_762 ();
 FILLCELL_X4 FILLER_153_766 ();
 FILLCELL_X8 FILLER_153_773 ();
 FILLCELL_X1 FILLER_153_791 ();
 FILLCELL_X1 FILLER_153_856 ();
 FILLCELL_X2 FILLER_153_859 ();
 FILLCELL_X1 FILLER_153_863 ();
 FILLCELL_X2 FILLER_153_884 ();
 FILLCELL_X4 FILLER_153_888 ();
 FILLCELL_X4 FILLER_153_899 ();
 FILLCELL_X4 FILLER_153_905 ();
 FILLCELL_X1 FILLER_153_929 ();
 FILLCELL_X8 FILLER_153_942 ();
 FILLCELL_X4 FILLER_153_950 ();
 FILLCELL_X2 FILLER_153_954 ();
 FILLCELL_X4 FILLER_153_974 ();
 FILLCELL_X8 FILLER_153_980 ();
 FILLCELL_X4 FILLER_153_988 ();
 FILLCELL_X1 FILLER_153_992 ();
 FILLCELL_X2 FILLER_153_996 ();
 FILLCELL_X1 FILLER_153_998 ();
 FILLCELL_X2 FILLER_153_1002 ();
 FILLCELL_X1 FILLER_153_1004 ();
 FILLCELL_X1 FILLER_153_1007 ();
 FILLCELL_X1 FILLER_153_1014 ();
 FILLCELL_X1 FILLER_153_1018 ();
 FILLCELL_X1 FILLER_153_1035 ();
 FILLCELL_X8 FILLER_153_1054 ();
 FILLCELL_X2 FILLER_153_1062 ();
 FILLCELL_X1 FILLER_153_1064 ();
 FILLCELL_X2 FILLER_153_1070 ();
 FILLCELL_X1 FILLER_153_1072 ();
 FILLCELL_X2 FILLER_153_1078 ();
 FILLCELL_X1 FILLER_153_1080 ();
 FILLCELL_X2 FILLER_153_1103 ();
 FILLCELL_X4 FILLER_153_1108 ();
 FILLCELL_X2 FILLER_153_1112 ();
 FILLCELL_X1 FILLER_153_1114 ();
 FILLCELL_X2 FILLER_153_1117 ();
 FILLCELL_X1 FILLER_153_1121 ();
 FILLCELL_X1 FILLER_153_1138 ();
 FILLCELL_X2 FILLER_153_1141 ();
 FILLCELL_X16 FILLER_153_1145 ();
 FILLCELL_X8 FILLER_153_1161 ();
 FILLCELL_X1 FILLER_153_1169 ();
 FILLCELL_X4 FILLER_153_1172 ();
 FILLCELL_X32 FILLER_153_1186 ();
 FILLCELL_X32 FILLER_153_1218 ();
 FILLCELL_X4 FILLER_153_1250 ();
 FILLCELL_X1 FILLER_153_1254 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X16 FILLER_154_321 ();
 FILLCELL_X8 FILLER_154_337 ();
 FILLCELL_X1 FILLER_154_345 ();
 FILLCELL_X8 FILLER_154_373 ();
 FILLCELL_X1 FILLER_154_381 ();
 FILLCELL_X8 FILLER_154_409 ();
 FILLCELL_X2 FILLER_154_417 ();
 FILLCELL_X1 FILLER_154_419 ();
 FILLCELL_X8 FILLER_154_447 ();
 FILLCELL_X1 FILLER_154_455 ();
 FILLCELL_X32 FILLER_154_483 ();
 FILLCELL_X32 FILLER_154_515 ();
 FILLCELL_X32 FILLER_154_547 ();
 FILLCELL_X32 FILLER_154_579 ();
 FILLCELL_X16 FILLER_154_611 ();
 FILLCELL_X4 FILLER_154_627 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X4 FILLER_154_696 ();
 FILLCELL_X2 FILLER_154_718 ();
 FILLCELL_X1 FILLER_154_720 ();
 FILLCELL_X2 FILLER_154_755 ();
 FILLCELL_X1 FILLER_154_757 ();
 FILLCELL_X1 FILLER_154_760 ();
 FILLCELL_X1 FILLER_154_763 ();
 FILLCELL_X1 FILLER_154_783 ();
 FILLCELL_X1 FILLER_154_800 ();
 FILLCELL_X8 FILLER_154_807 ();
 FILLCELL_X2 FILLER_154_815 ();
 FILLCELL_X4 FILLER_154_819 ();
 FILLCELL_X1 FILLER_154_823 ();
 FILLCELL_X2 FILLER_154_828 ();
 FILLCELL_X1 FILLER_154_830 ();
 FILLCELL_X8 FILLER_154_834 ();
 FILLCELL_X2 FILLER_154_842 ();
 FILLCELL_X16 FILLER_154_846 ();
 FILLCELL_X1 FILLER_154_862 ();
 FILLCELL_X1 FILLER_154_881 ();
 FILLCELL_X2 FILLER_154_884 ();
 FILLCELL_X1 FILLER_154_886 ();
 FILLCELL_X4 FILLER_154_931 ();
 FILLCELL_X4 FILLER_154_969 ();
 FILLCELL_X2 FILLER_154_973 ();
 FILLCELL_X4 FILLER_154_977 ();
 FILLCELL_X1 FILLER_154_984 ();
 FILLCELL_X2 FILLER_154_1017 ();
 FILLCELL_X4 FILLER_154_1024 ();
 FILLCELL_X1 FILLER_154_1028 ();
 FILLCELL_X8 FILLER_154_1031 ();
 FILLCELL_X1 FILLER_154_1096 ();
 FILLCELL_X1 FILLER_154_1113 ();
 FILLCELL_X1 FILLER_154_1130 ();
 FILLCELL_X1 FILLER_154_1147 ();
 FILLCELL_X2 FILLER_154_1160 ();
 FILLCELL_X1 FILLER_154_1162 ();
 FILLCELL_X4 FILLER_154_1167 ();
 FILLCELL_X2 FILLER_154_1171 ();
 FILLCELL_X1 FILLER_154_1180 ();
 FILLCELL_X32 FILLER_154_1191 ();
 FILLCELL_X32 FILLER_154_1223 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X16 FILLER_155_673 ();
 FILLCELL_X8 FILLER_155_689 ();
 FILLCELL_X4 FILLER_155_697 ();
 FILLCELL_X2 FILLER_155_701 ();
 FILLCELL_X1 FILLER_155_703 ();
 FILLCELL_X8 FILLER_155_738 ();
 FILLCELL_X2 FILLER_155_746 ();
 FILLCELL_X4 FILLER_155_750 ();
 FILLCELL_X2 FILLER_155_754 ();
 FILLCELL_X1 FILLER_155_756 ();
 FILLCELL_X8 FILLER_155_759 ();
 FILLCELL_X2 FILLER_155_783 ();
 FILLCELL_X4 FILLER_155_787 ();
 FILLCELL_X1 FILLER_155_791 ();
 FILLCELL_X2 FILLER_155_816 ();
 FILLCELL_X16 FILLER_155_836 ();
 FILLCELL_X1 FILLER_155_852 ();
 FILLCELL_X2 FILLER_155_869 ();
 FILLCELL_X1 FILLER_155_871 ();
 FILLCELL_X16 FILLER_155_906 ();
 FILLCELL_X1 FILLER_155_922 ();
 FILLCELL_X2 FILLER_155_925 ();
 FILLCELL_X2 FILLER_155_947 ();
 FILLCELL_X1 FILLER_155_949 ();
 FILLCELL_X8 FILLER_155_952 ();
 FILLCELL_X4 FILLER_155_960 ();
 FILLCELL_X2 FILLER_155_964 ();
 FILLCELL_X1 FILLER_155_966 ();
 FILLCELL_X2 FILLER_155_969 ();
 FILLCELL_X8 FILLER_155_990 ();
 FILLCELL_X2 FILLER_155_998 ();
 FILLCELL_X1 FILLER_155_1000 ();
 FILLCELL_X1 FILLER_155_1004 ();
 FILLCELL_X8 FILLER_155_1007 ();
 FILLCELL_X2 FILLER_155_1015 ();
 FILLCELL_X1 FILLER_155_1040 ();
 FILLCELL_X2 FILLER_155_1057 ();
 FILLCELL_X1 FILLER_155_1062 ();
 FILLCELL_X2 FILLER_155_1069 ();
 FILLCELL_X1 FILLER_155_1074 ();
 FILLCELL_X4 FILLER_155_1101 ();
 FILLCELL_X1 FILLER_155_1105 ();
 FILLCELL_X2 FILLER_155_1109 ();
 FILLCELL_X1 FILLER_155_1111 ();
 FILLCELL_X8 FILLER_155_1115 ();
 FILLCELL_X4 FILLER_155_1123 ();
 FILLCELL_X2 FILLER_155_1127 ();
 FILLCELL_X8 FILLER_155_1139 ();
 FILLCELL_X2 FILLER_155_1147 ();
 FILLCELL_X1 FILLER_155_1149 ();
 FILLCELL_X4 FILLER_155_1166 ();
 FILLCELL_X2 FILLER_155_1170 ();
 FILLCELL_X32 FILLER_155_1188 ();
 FILLCELL_X32 FILLER_155_1220 ();
 FILLCELL_X2 FILLER_155_1252 ();
 FILLCELL_X1 FILLER_155_1254 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X8 FILLER_156_696 ();
 FILLCELL_X2 FILLER_156_704 ();
 FILLCELL_X1 FILLER_156_706 ();
 FILLCELL_X2 FILLER_156_715 ();
 FILLCELL_X1 FILLER_156_717 ();
 FILLCELL_X8 FILLER_156_800 ();
 FILLCELL_X4 FILLER_156_808 ();
 FILLCELL_X2 FILLER_156_812 ();
 FILLCELL_X1 FILLER_156_814 ();
 FILLCELL_X2 FILLER_156_831 ();
 FILLCELL_X1 FILLER_156_833 ();
 FILLCELL_X16 FILLER_156_866 ();
 FILLCELL_X4 FILLER_156_882 ();
 FILLCELL_X2 FILLER_156_886 ();
 FILLCELL_X4 FILLER_156_891 ();
 FILLCELL_X2 FILLER_156_895 ();
 FILLCELL_X4 FILLER_156_913 ();
 FILLCELL_X2 FILLER_156_917 ();
 FILLCELL_X4 FILLER_156_935 ();
 FILLCELL_X2 FILLER_156_939 ();
 FILLCELL_X1 FILLER_156_960 ();
 FILLCELL_X8 FILLER_156_964 ();
 FILLCELL_X2 FILLER_156_1019 ();
 FILLCELL_X1 FILLER_156_1024 ();
 FILLCELL_X2 FILLER_156_1060 ();
 FILLCELL_X1 FILLER_156_1062 ();
 FILLCELL_X8 FILLER_156_1094 ();
 FILLCELL_X1 FILLER_156_1102 ();
 FILLCELL_X32 FILLER_156_1124 ();
 FILLCELL_X8 FILLER_156_1156 ();
 FILLCELL_X4 FILLER_156_1164 ();
 FILLCELL_X1 FILLER_156_1168 ();
 FILLCELL_X32 FILLER_156_1186 ();
 FILLCELL_X32 FILLER_156_1218 ();
 FILLCELL_X4 FILLER_156_1250 ();
 FILLCELL_X1 FILLER_156_1254 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X4 FILLER_157_737 ();
 FILLCELL_X4 FILLER_157_773 ();
 FILLCELL_X2 FILLER_157_777 ();
 FILLCELL_X4 FILLER_157_843 ();
 FILLCELL_X2 FILLER_157_847 ();
 FILLCELL_X2 FILLER_157_857 ();
 FILLCELL_X1 FILLER_157_859 ();
 FILLCELL_X8 FILLER_157_878 ();
 FILLCELL_X4 FILLER_157_886 ();
 FILLCELL_X4 FILLER_157_892 ();
 FILLCELL_X2 FILLER_157_896 ();
 FILLCELL_X2 FILLER_157_900 ();
 FILLCELL_X8 FILLER_157_904 ();
 FILLCELL_X2 FILLER_157_912 ();
 FILLCELL_X2 FILLER_157_917 ();
 FILLCELL_X1 FILLER_157_919 ();
 FILLCELL_X8 FILLER_157_923 ();
 FILLCELL_X2 FILLER_157_931 ();
 FILLCELL_X1 FILLER_157_933 ();
 FILLCELL_X4 FILLER_157_940 ();
 FILLCELL_X2 FILLER_157_944 ();
 FILLCELL_X4 FILLER_157_948 ();
 FILLCELL_X1 FILLER_157_1000 ();
 FILLCELL_X2 FILLER_157_1033 ();
 FILLCELL_X4 FILLER_157_1075 ();
 FILLCELL_X1 FILLER_157_1079 ();
 FILLCELL_X4 FILLER_157_1101 ();
 FILLCELL_X1 FILLER_157_1105 ();
 FILLCELL_X2 FILLER_157_1114 ();
 FILLCELL_X1 FILLER_157_1132 ();
 FILLCELL_X1 FILLER_157_1165 ();
 FILLCELL_X32 FILLER_157_1189 ();
 FILLCELL_X32 FILLER_157_1221 ();
 FILLCELL_X2 FILLER_157_1253 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X16 FILLER_158_696 ();
 FILLCELL_X2 FILLER_158_712 ();
 FILLCELL_X16 FILLER_158_748 ();
 FILLCELL_X4 FILLER_158_764 ();
 FILLCELL_X16 FILLER_158_784 ();
 FILLCELL_X2 FILLER_158_819 ();
 FILLCELL_X4 FILLER_158_835 ();
 FILLCELL_X2 FILLER_158_848 ();
 FILLCELL_X2 FILLER_158_852 ();
 FILLCELL_X1 FILLER_158_854 ();
 FILLCELL_X1 FILLER_158_857 ();
 FILLCELL_X1 FILLER_158_874 ();
 FILLCELL_X1 FILLER_158_891 ();
 FILLCELL_X2 FILLER_158_943 ();
 FILLCELL_X1 FILLER_158_945 ();
 FILLCELL_X4 FILLER_158_949 ();
 FILLCELL_X1 FILLER_158_976 ();
 FILLCELL_X4 FILLER_158_993 ();
 FILLCELL_X8 FILLER_158_1013 ();
 FILLCELL_X2 FILLER_158_1021 ();
 FILLCELL_X1 FILLER_158_1023 ();
 FILLCELL_X2 FILLER_158_1056 ();
 FILLCELL_X1 FILLER_158_1058 ();
 FILLCELL_X1 FILLER_158_1078 ();
 FILLCELL_X4 FILLER_158_1098 ();
 FILLCELL_X2 FILLER_158_1121 ();
 FILLCELL_X4 FILLER_158_1135 ();
 FILLCELL_X1 FILLER_158_1139 ();
 FILLCELL_X1 FILLER_158_1156 ();
 FILLCELL_X32 FILLER_158_1179 ();
 FILLCELL_X32 FILLER_158_1211 ();
 FILLCELL_X8 FILLER_158_1243 ();
 FILLCELL_X4 FILLER_158_1251 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X16 FILLER_159_705 ();
 FILLCELL_X2 FILLER_159_721 ();
 FILLCELL_X8 FILLER_159_725 ();
 FILLCELL_X4 FILLER_159_733 ();
 FILLCELL_X2 FILLER_159_737 ();
 FILLCELL_X8 FILLER_159_741 ();
 FILLCELL_X4 FILLER_159_765 ();
 FILLCELL_X2 FILLER_159_769 ();
 FILLCELL_X1 FILLER_159_771 ();
 FILLCELL_X4 FILLER_159_827 ();
 FILLCELL_X2 FILLER_159_863 ();
 FILLCELL_X8 FILLER_159_901 ();
 FILLCELL_X1 FILLER_159_913 ();
 FILLCELL_X2 FILLER_159_930 ();
 FILLCELL_X4 FILLER_159_964 ();
 FILLCELL_X1 FILLER_159_968 ();
 FILLCELL_X1 FILLER_159_972 ();
 FILLCELL_X4 FILLER_159_976 ();
 FILLCELL_X8 FILLER_159_1028 ();
 FILLCELL_X4 FILLER_159_1036 ();
 FILLCELL_X2 FILLER_159_1040 ();
 FILLCELL_X8 FILLER_159_1116 ();
 FILLCELL_X1 FILLER_159_1124 ();
 FILLCELL_X1 FILLER_159_1145 ();
 FILLCELL_X2 FILLER_159_1150 ();
 FILLCELL_X1 FILLER_159_1152 ();
 FILLCELL_X2 FILLER_159_1155 ();
 FILLCELL_X2 FILLER_159_1159 ();
 FILLCELL_X1 FILLER_159_1161 ();
 FILLCELL_X32 FILLER_159_1178 ();
 FILLCELL_X32 FILLER_159_1210 ();
 FILLCELL_X8 FILLER_159_1242 ();
 FILLCELL_X4 FILLER_159_1250 ();
 FILLCELL_X1 FILLER_159_1254 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X16 FILLER_160_744 ();
 FILLCELL_X1 FILLER_160_783 ();
 FILLCELL_X16 FILLER_160_803 ();
 FILLCELL_X8 FILLER_160_819 ();
 FILLCELL_X1 FILLER_160_827 ();
 FILLCELL_X8 FILLER_160_833 ();
 FILLCELL_X8 FILLER_160_852 ();
 FILLCELL_X2 FILLER_160_860 ();
 FILLCELL_X8 FILLER_160_868 ();
 FILLCELL_X2 FILLER_160_894 ();
 FILLCELL_X4 FILLER_160_919 ();
 FILLCELL_X1 FILLER_160_923 ();
 FILLCELL_X2 FILLER_160_940 ();
 FILLCELL_X1 FILLER_160_942 ();
 FILLCELL_X32 FILLER_160_946 ();
 FILLCELL_X32 FILLER_160_978 ();
 FILLCELL_X8 FILLER_160_1010 ();
 FILLCELL_X2 FILLER_160_1018 ();
 FILLCELL_X2 FILLER_160_1036 ();
 FILLCELL_X1 FILLER_160_1038 ();
 FILLCELL_X4 FILLER_160_1055 ();
 FILLCELL_X8 FILLER_160_1079 ();
 FILLCELL_X2 FILLER_160_1087 ();
 FILLCELL_X1 FILLER_160_1089 ();
 FILLCELL_X2 FILLER_160_1108 ();
 FILLCELL_X1 FILLER_160_1110 ();
 FILLCELL_X8 FILLER_160_1113 ();
 FILLCELL_X2 FILLER_160_1121 ();
 FILLCELL_X1 FILLER_160_1123 ();
 FILLCELL_X1 FILLER_160_1140 ();
 FILLCELL_X1 FILLER_160_1143 ();
 FILLCELL_X2 FILLER_160_1165 ();
 FILLCELL_X32 FILLER_160_1177 ();
 FILLCELL_X32 FILLER_160_1209 ();
 FILLCELL_X8 FILLER_160_1241 ();
 FILLCELL_X4 FILLER_160_1249 ();
 FILLCELL_X2 FILLER_160_1253 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X4 FILLER_161_737 ();
 FILLCELL_X1 FILLER_161_741 ();
 FILLCELL_X1 FILLER_161_760 ();
 FILLCELL_X1 FILLER_161_775 ();
 FILLCELL_X2 FILLER_161_779 ();
 FILLCELL_X1 FILLER_161_784 ();
 FILLCELL_X1 FILLER_161_801 ();
 FILLCELL_X2 FILLER_161_805 ();
 FILLCELL_X1 FILLER_161_807 ();
 FILLCELL_X8 FILLER_161_811 ();
 FILLCELL_X4 FILLER_161_819 ();
 FILLCELL_X4 FILLER_161_832 ();
 FILLCELL_X16 FILLER_161_871 ();
 FILLCELL_X8 FILLER_161_887 ();
 FILLCELL_X1 FILLER_161_895 ();
 FILLCELL_X8 FILLER_161_899 ();
 FILLCELL_X4 FILLER_161_907 ();
 FILLCELL_X2 FILLER_161_911 ();
 FILLCELL_X2 FILLER_161_929 ();
 FILLCELL_X1 FILLER_161_931 ();
 FILLCELL_X16 FILLER_161_948 ();
 FILLCELL_X2 FILLER_161_964 ();
 FILLCELL_X1 FILLER_161_966 ();
 FILLCELL_X4 FILLER_161_983 ();
 FILLCELL_X1 FILLER_161_987 ();
 FILLCELL_X4 FILLER_161_1004 ();
 FILLCELL_X2 FILLER_161_1008 ();
 FILLCELL_X4 FILLER_161_1016 ();
 FILLCELL_X2 FILLER_161_1020 ();
 FILLCELL_X8 FILLER_161_1034 ();
 FILLCELL_X4 FILLER_161_1084 ();
 FILLCELL_X1 FILLER_161_1088 ();
 FILLCELL_X4 FILLER_161_1157 ();
 FILLCELL_X2 FILLER_161_1161 ();
 FILLCELL_X32 FILLER_161_1167 ();
 FILLCELL_X32 FILLER_161_1199 ();
 FILLCELL_X16 FILLER_161_1231 ();
 FILLCELL_X8 FILLER_161_1247 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X16 FILLER_162_728 ();
 FILLCELL_X8 FILLER_162_744 ();
 FILLCELL_X4 FILLER_162_752 ();
 FILLCELL_X2 FILLER_162_756 ();
 FILLCELL_X1 FILLER_162_758 ();
 FILLCELL_X8 FILLER_162_766 ();
 FILLCELL_X4 FILLER_162_774 ();
 FILLCELL_X2 FILLER_162_778 ();
 FILLCELL_X1 FILLER_162_780 ();
 FILLCELL_X1 FILLER_162_835 ();
 FILLCELL_X4 FILLER_162_839 ();
 FILLCELL_X1 FILLER_162_846 ();
 FILLCELL_X2 FILLER_162_863 ();
 FILLCELL_X2 FILLER_162_868 ();
 FILLCELL_X2 FILLER_162_873 ();
 FILLCELL_X1 FILLER_162_875 ();
 FILLCELL_X4 FILLER_162_879 ();
 FILLCELL_X1 FILLER_162_883 ();
 FILLCELL_X8 FILLER_162_887 ();
 FILLCELL_X2 FILLER_162_895 ();
 FILLCELL_X2 FILLER_162_900 ();
 FILLCELL_X1 FILLER_162_902 ();
 FILLCELL_X2 FILLER_162_926 ();
 FILLCELL_X8 FILLER_162_992 ();
 FILLCELL_X2 FILLER_162_1000 ();
 FILLCELL_X2 FILLER_162_1037 ();
 FILLCELL_X1 FILLER_162_1039 ();
 FILLCELL_X8 FILLER_162_1042 ();
 FILLCELL_X2 FILLER_162_1050 ();
 FILLCELL_X1 FILLER_162_1052 ();
 FILLCELL_X2 FILLER_162_1070 ();
 FILLCELL_X4 FILLER_162_1074 ();
 FILLCELL_X2 FILLER_162_1078 ();
 FILLCELL_X8 FILLER_162_1096 ();
 FILLCELL_X1 FILLER_162_1104 ();
 FILLCELL_X1 FILLER_162_1111 ();
 FILLCELL_X4 FILLER_162_1115 ();
 FILLCELL_X2 FILLER_162_1119 ();
 FILLCELL_X1 FILLER_162_1123 ();
 FILLCELL_X1 FILLER_162_1140 ();
 FILLCELL_X32 FILLER_162_1162 ();
 FILLCELL_X32 FILLER_162_1194 ();
 FILLCELL_X16 FILLER_162_1226 ();
 FILLCELL_X8 FILLER_162_1242 ();
 FILLCELL_X4 FILLER_162_1250 ();
 FILLCELL_X1 FILLER_162_1254 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X16 FILLER_163_737 ();
 FILLCELL_X8 FILLER_163_753 ();
 FILLCELL_X4 FILLER_163_761 ();
 FILLCELL_X2 FILLER_163_765 ();
 FILLCELL_X1 FILLER_163_767 ();
 FILLCELL_X2 FILLER_163_771 ();
 FILLCELL_X2 FILLER_163_777 ();
 FILLCELL_X8 FILLER_163_782 ();
 FILLCELL_X4 FILLER_163_790 ();
 FILLCELL_X2 FILLER_163_794 ();
 FILLCELL_X8 FILLER_163_954 ();
 FILLCELL_X2 FILLER_163_962 ();
 FILLCELL_X4 FILLER_163_969 ();
 FILLCELL_X2 FILLER_163_973 ();
 FILLCELL_X2 FILLER_163_978 ();
 FILLCELL_X4 FILLER_163_996 ();
 FILLCELL_X2 FILLER_163_1000 ();
 FILLCELL_X2 FILLER_163_1021 ();
 FILLCELL_X2 FILLER_163_1041 ();
 FILLCELL_X1 FILLER_163_1056 ();
 FILLCELL_X4 FILLER_163_1061 ();
 FILLCELL_X4 FILLER_163_1075 ();
 FILLCELL_X2 FILLER_163_1092 ();
 FILLCELL_X1 FILLER_163_1094 ();
 FILLCELL_X2 FILLER_163_1098 ();
 FILLCELL_X1 FILLER_163_1100 ();
 FILLCELL_X2 FILLER_163_1120 ();
 FILLCELL_X8 FILLER_163_1124 ();
 FILLCELL_X4 FILLER_163_1142 ();
 FILLCELL_X2 FILLER_163_1146 ();
 FILLCELL_X1 FILLER_163_1148 ();
 FILLCELL_X32 FILLER_163_1151 ();
 FILLCELL_X32 FILLER_163_1183 ();
 FILLCELL_X32 FILLER_163_1215 ();
 FILLCELL_X8 FILLER_163_1247 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X4 FILLER_164_760 ();
 FILLCELL_X2 FILLER_164_764 ();
 FILLCELL_X1 FILLER_164_766 ();
 FILLCELL_X8 FILLER_164_785 ();
 FILLCELL_X8 FILLER_164_796 ();
 FILLCELL_X4 FILLER_164_812 ();
 FILLCELL_X1 FILLER_164_816 ();
 FILLCELL_X4 FILLER_164_833 ();
 FILLCELL_X2 FILLER_164_837 ();
 FILLCELL_X1 FILLER_164_839 ();
 FILLCELL_X8 FILLER_164_843 ();
 FILLCELL_X4 FILLER_164_861 ();
 FILLCELL_X2 FILLER_164_865 ();
 FILLCELL_X8 FILLER_164_873 ();
 FILLCELL_X4 FILLER_164_881 ();
 FILLCELL_X8 FILLER_164_888 ();
 FILLCELL_X1 FILLER_164_901 ();
 FILLCELL_X4 FILLER_164_904 ();
 FILLCELL_X1 FILLER_164_908 ();
 FILLCELL_X2 FILLER_164_912 ();
 FILLCELL_X8 FILLER_164_920 ();
 FILLCELL_X4 FILLER_164_928 ();
 FILLCELL_X4 FILLER_164_967 ();
 FILLCELL_X1 FILLER_164_971 ();
 FILLCELL_X2 FILLER_164_978 ();
 FILLCELL_X1 FILLER_164_1028 ();
 FILLCELL_X2 FILLER_164_1063 ();
 FILLCELL_X1 FILLER_164_1065 ();
 FILLCELL_X4 FILLER_164_1085 ();
 FILLCELL_X2 FILLER_164_1089 ();
 FILLCELL_X4 FILLER_164_1094 ();
 FILLCELL_X1 FILLER_164_1098 ();
 FILLCELL_X2 FILLER_164_1105 ();
 FILLCELL_X1 FILLER_164_1107 ();
 FILLCELL_X8 FILLER_164_1111 ();
 FILLCELL_X1 FILLER_164_1121 ();
 FILLCELL_X32 FILLER_164_1142 ();
 FILLCELL_X32 FILLER_164_1174 ();
 FILLCELL_X32 FILLER_164_1206 ();
 FILLCELL_X16 FILLER_164_1238 ();
 FILLCELL_X1 FILLER_164_1254 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X8 FILLER_165_804 ();
 FILLCELL_X4 FILLER_165_812 ();
 FILLCELL_X2 FILLER_165_816 ();
 FILLCELL_X1 FILLER_165_818 ();
 FILLCELL_X8 FILLER_165_822 ();
 FILLCELL_X2 FILLER_165_830 ();
 FILLCELL_X1 FILLER_165_832 ();
 FILLCELL_X2 FILLER_165_849 ();
 FILLCELL_X1 FILLER_165_851 ();
 FILLCELL_X4 FILLER_165_886 ();
 FILLCELL_X2 FILLER_165_890 ();
 FILLCELL_X4 FILLER_165_941 ();
 FILLCELL_X4 FILLER_165_947 ();
 FILLCELL_X2 FILLER_165_951 ();
 FILLCELL_X4 FILLER_165_959 ();
 FILLCELL_X2 FILLER_165_963 ();
 FILLCELL_X1 FILLER_165_965 ();
 FILLCELL_X4 FILLER_165_984 ();
 FILLCELL_X2 FILLER_165_988 ();
 FILLCELL_X1 FILLER_165_992 ();
 FILLCELL_X2 FILLER_165_996 ();
 FILLCELL_X1 FILLER_165_1001 ();
 FILLCELL_X4 FILLER_165_1005 ();
 FILLCELL_X1 FILLER_165_1009 ();
 FILLCELL_X4 FILLER_165_1012 ();
 FILLCELL_X1 FILLER_165_1016 ();
 FILLCELL_X2 FILLER_165_1020 ();
 FILLCELL_X2 FILLER_165_1024 ();
 FILLCELL_X2 FILLER_165_1029 ();
 FILLCELL_X4 FILLER_165_1037 ();
 FILLCELL_X2 FILLER_165_1041 ();
 FILLCELL_X1 FILLER_165_1043 ();
 FILLCELL_X2 FILLER_165_1050 ();
 FILLCELL_X1 FILLER_165_1055 ();
 FILLCELL_X1 FILLER_165_1074 ();
 FILLCELL_X1 FILLER_165_1091 ();
 FILLCELL_X1 FILLER_165_1095 ();
 FILLCELL_X2 FILLER_165_1106 ();
 FILLCELL_X2 FILLER_165_1127 ();
 FILLCELL_X1 FILLER_165_1129 ();
 FILLCELL_X1 FILLER_165_1132 ();
 FILLCELL_X32 FILLER_165_1143 ();
 FILLCELL_X32 FILLER_165_1175 ();
 FILLCELL_X32 FILLER_165_1207 ();
 FILLCELL_X16 FILLER_165_1239 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X2 FILLER_166_792 ();
 FILLCELL_X16 FILLER_166_842 ();
 FILLCELL_X8 FILLER_166_858 ();
 FILLCELL_X2 FILLER_166_866 ();
 FILLCELL_X1 FILLER_166_868 ();
 FILLCELL_X4 FILLER_166_906 ();
 FILLCELL_X4 FILLER_166_916 ();
 FILLCELL_X4 FILLER_166_922 ();
 FILLCELL_X2 FILLER_166_926 ();
 FILLCELL_X8 FILLER_166_934 ();
 FILLCELL_X1 FILLER_166_942 ();
 FILLCELL_X2 FILLER_166_945 ();
 FILLCELL_X4 FILLER_166_963 ();
 FILLCELL_X2 FILLER_166_967 ();
 FILLCELL_X1 FILLER_166_969 ();
 FILLCELL_X1 FILLER_166_972 ();
 FILLCELL_X8 FILLER_166_976 ();
 FILLCELL_X1 FILLER_166_984 ();
 FILLCELL_X8 FILLER_166_1010 ();
 FILLCELL_X2 FILLER_166_1018 ();
 FILLCELL_X1 FILLER_166_1020 ();
 FILLCELL_X2 FILLER_166_1037 ();
 FILLCELL_X16 FILLER_166_1058 ();
 FILLCELL_X2 FILLER_166_1074 ();
 FILLCELL_X1 FILLER_166_1076 ();
 FILLCELL_X2 FILLER_166_1079 ();
 FILLCELL_X1 FILLER_166_1081 ();
 FILLCELL_X8 FILLER_166_1087 ();
 FILLCELL_X4 FILLER_166_1095 ();
 FILLCELL_X2 FILLER_166_1099 ();
 FILLCELL_X1 FILLER_166_1101 ();
 FILLCELL_X2 FILLER_166_1105 ();
 FILLCELL_X1 FILLER_166_1107 ();
 FILLCELL_X4 FILLER_166_1111 ();
 FILLCELL_X1 FILLER_166_1115 ();
 FILLCELL_X4 FILLER_166_1118 ();
 FILLCELL_X2 FILLER_166_1122 ();
 FILLCELL_X1 FILLER_166_1124 ();
 FILLCELL_X32 FILLER_166_1137 ();
 FILLCELL_X32 FILLER_166_1169 ();
 FILLCELL_X32 FILLER_166_1201 ();
 FILLCELL_X16 FILLER_166_1233 ();
 FILLCELL_X4 FILLER_166_1249 ();
 FILLCELL_X2 FILLER_166_1253 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X2 FILLER_167_801 ();
 FILLCELL_X8 FILLER_167_806 ();
 FILLCELL_X1 FILLER_167_836 ();
 FILLCELL_X2 FILLER_167_840 ();
 FILLCELL_X4 FILLER_167_877 ();
 FILLCELL_X2 FILLER_167_881 ();
 FILLCELL_X1 FILLER_167_883 ();
 FILLCELL_X1 FILLER_167_887 ();
 FILLCELL_X4 FILLER_167_891 ();
 FILLCELL_X2 FILLER_167_911 ();
 FILLCELL_X1 FILLER_167_916 ();
 FILLCELL_X2 FILLER_167_920 ();
 FILLCELL_X1 FILLER_167_938 ();
 FILLCELL_X1 FILLER_167_961 ();
 FILLCELL_X8 FILLER_167_997 ();
 FILLCELL_X4 FILLER_167_1005 ();
 FILLCELL_X2 FILLER_167_1009 ();
 FILLCELL_X4 FILLER_167_1014 ();
 FILLCELL_X8 FILLER_167_1020 ();
 FILLCELL_X8 FILLER_167_1034 ();
 FILLCELL_X16 FILLER_167_1044 ();
 FILLCELL_X4 FILLER_167_1066 ();
 FILLCELL_X1 FILLER_167_1070 ();
 FILLCELL_X2 FILLER_167_1087 ();
 FILLCELL_X4 FILLER_167_1095 ();
 FILLCELL_X2 FILLER_167_1099 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X4 FILLER_167_1249 ();
 FILLCELL_X2 FILLER_167_1253 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X1 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_636 ();
 FILLCELL_X32 FILLER_168_668 ();
 FILLCELL_X32 FILLER_168_700 ();
 FILLCELL_X32 FILLER_168_732 ();
 FILLCELL_X32 FILLER_168_764 ();
 FILLCELL_X32 FILLER_168_796 ();
 FILLCELL_X8 FILLER_168_828 ();
 FILLCELL_X2 FILLER_168_852 ();
 FILLCELL_X4 FILLER_168_857 ();
 FILLCELL_X2 FILLER_168_861 ();
 FILLCELL_X2 FILLER_168_879 ();
 FILLCELL_X2 FILLER_168_932 ();
 FILLCELL_X1 FILLER_168_934 ();
 FILLCELL_X1 FILLER_168_954 ();
 FILLCELL_X8 FILLER_168_974 ();
 FILLCELL_X2 FILLER_168_982 ();
 FILLCELL_X32 FILLER_168_1121 ();
 FILLCELL_X32 FILLER_168_1153 ();
 FILLCELL_X32 FILLER_168_1185 ();
 FILLCELL_X32 FILLER_168_1217 ();
 FILLCELL_X4 FILLER_168_1249 ();
 FILLCELL_X2 FILLER_168_1253 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X2 FILLER_169_577 ();
 FILLCELL_X1 FILLER_169_579 ();
 FILLCELL_X2 FILLER_169_583 ();
 FILLCELL_X1 FILLER_169_585 ();
 FILLCELL_X2 FILLER_169_598 ();
 FILLCELL_X1 FILLER_169_600 ();
 FILLCELL_X2 FILLER_169_625 ();
 FILLCELL_X1 FILLER_169_627 ();
 FILLCELL_X4 FILLER_169_632 ();
 FILLCELL_X1 FILLER_169_636 ();
 FILLCELL_X32 FILLER_169_643 ();
 FILLCELL_X32 FILLER_169_675 ();
 FILLCELL_X32 FILLER_169_707 ();
 FILLCELL_X32 FILLER_169_739 ();
 FILLCELL_X32 FILLER_169_771 ();
 FILLCELL_X32 FILLER_169_803 ();
 FILLCELL_X32 FILLER_169_835 ();
 FILLCELL_X16 FILLER_169_870 ();
 FILLCELL_X2 FILLER_169_886 ();
 FILLCELL_X8 FILLER_169_891 ();
 FILLCELL_X2 FILLER_169_899 ();
 FILLCELL_X2 FILLER_169_914 ();
 FILLCELL_X8 FILLER_169_932 ();
 FILLCELL_X1 FILLER_169_940 ();
 FILLCELL_X16 FILLER_169_944 ();
 FILLCELL_X2 FILLER_169_960 ();
 FILLCELL_X1 FILLER_169_962 ();
 FILLCELL_X16 FILLER_169_966 ();
 FILLCELL_X8 FILLER_169_982 ();
 FILLCELL_X4 FILLER_169_990 ();
 FILLCELL_X2 FILLER_169_994 ();
 FILLCELL_X16 FILLER_169_1005 ();
 FILLCELL_X4 FILLER_169_1021 ();
 FILLCELL_X1 FILLER_169_1025 ();
 FILLCELL_X16 FILLER_169_1032 ();
 FILLCELL_X4 FILLER_169_1048 ();
 FILLCELL_X1 FILLER_169_1052 ();
 FILLCELL_X4 FILLER_169_1055 ();
 FILLCELL_X2 FILLER_169_1059 ();
 FILLCELL_X8 FILLER_169_1064 ();
 FILLCELL_X2 FILLER_169_1072 ();
 FILLCELL_X1 FILLER_169_1074 ();
 FILLCELL_X4 FILLER_169_1087 ();
 FILLCELL_X2 FILLER_169_1091 ();
 FILLCELL_X1 FILLER_169_1093 ();
 FILLCELL_X32 FILLER_169_1097 ();
 FILLCELL_X32 FILLER_169_1129 ();
 FILLCELL_X32 FILLER_169_1161 ();
 FILLCELL_X32 FILLER_169_1193 ();
 FILLCELL_X16 FILLER_169_1225 ();
 FILLCELL_X8 FILLER_169_1241 ();
 FILLCELL_X4 FILLER_169_1249 ();
 FILLCELL_X2 FILLER_169_1253 ();
endmodule
