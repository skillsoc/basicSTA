//
// Conformal-LEC: Version 07.20-d165 (10-Mar-2008)
//
module rom_512x16A(Q, CLK, CEN, A);
// dont_use
input  CLK, CEN;
input   [8:0] A;
output  [15:0] Q;
  // module is bboxed.
endmodule

