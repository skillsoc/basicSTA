//
// Conformal-LEC: Version 07.20-d165 (10-Mar-2008)
//
module ram_256x16A(Q, CLK, CEN, WEN, A, D);
// dont_use
input  CLK, CEN, WEN;
input   [7:0] A;
input   [15:0] D;
output  [15:0] Q;
  // module is bboxed.
endmodule

