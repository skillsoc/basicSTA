VERSION   5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
   DATABASE MICRONS 2000 ;
END UNITS

MACRO pllclk
  CLASS BLOCK ;
  ORIGIN 0.06 0 ;
  SIZE 150.06 BY 273.59 ;
  SYMMETRY X Y R90 ;

  PIN refclk
  DIRECTION INPUT ;
     PORT
      LAYER M1 ;
      RECT 0 160.23 0.3 160.61 ;
     END
  END refclk

  PIN clk1x
  DIRECTION OUTPUT ;
     PORT
      LAYER M2 ;
      RECT 63.72 226.08 64.32 226.68 ;
     END
  END clk1x

  PIN clk2x
  DIRECTION OUTPUT ;
     PORT
      LAYER M2 ;
      RECT 63.72 244.56 64.32 245.16 ;
     END
  END clk2x

  PIN ibias
  DIRECTION INPUT ;
     PORT
      LAYER M2 ;
      RECT 0 179.9 0.6 180.5 ;
     END
  END ibias

  PIN reset
  DIRECTION INPUT ;
     PORT
      LAYER M2 ;
      RECT 0 182.54 0.6 183.14 ;
     END
  END reset

  PIN vcom
  DIRECTION OUTPUT ;
     PORT
      LAYER M2 ;
      RECT 0 174.62 0.6 175.22 ;
     END
  END vcom

  PIN vcop
  DIRECTION OUTPUT ;
     PORT
      LAYER M2 ;
      RECT 0 177.26 0.6 177.86 ;
     END
  END vcop

  PIN agnd!
  DIRECTION INOUT ;
  USE GROUND ;
     PORT
      LAYER M3 ;
      RECT 0 4.78 132.28 9.78 ;
      RECT 0 4.77 0.6 9.78 ;
     END
     PORT
      LAYER M3 ;
      RECT 0 168.46 132.28 173.46 ;
     END
  END agnd!

  PIN avdd!
  DIRECTION INOUT ;
  USE POWER ;
     PORT
      LAYER M3 ;
      RECT 0 11.37 0.6 16.38 ;
      RECT 0 11.38 132.28 16.38 ;
     END
     PORT
      LAYER M3 ;
      RECT 0 161.85 0.59 166.86 ;
      RECT -0.01 161.86 132.28 166.85 ;
      RECT -0.01 161.85 0.59 166.85 ;
      RECT 0 161.86 132.28 166.86 ;
     END
  END avdd!
  OBS
      LAYER OVERLAP ;
      POLYGON 150 173.46 68.64 173.46 68.64 217.03 64.32 217.03 64.32 273.59 0 273.59 0 0 150 0 ;
#  POLYGON 150 173.46 68.64 173.46 68.64 217.03 64.32 217.03 64.32 273.59 10.49 273.59 10.49 206.26 0 206.26 0 0 150 0 ;
      LAYER M1 ;
      POLYGON 149.885 173.345 68.525 173.345 68.525 216.915 64.205 216.915 64.205 273.475 10.605 273.475 10.605 206.145 0.115 206.145 0.115 160.84 0.53 160.84 0.53 160
         0.115 160 0.115 159.21 0 159.21 0 158.91 0.115 158.91 0.115 0.115 149.885 0.115 ;
      LAYER M2 ;
      POLYGON 149.86 173.32 68.5 173.32 68.5 216.89 64.18 216.89 64.18 225.8 63.44 225.8 63.44 226.96 64.18 226.96 64.18 244.28 63.44 244.28 63.44 245.44
         64.18 245.44 64.18 263.04 64.32 263.04 64.32 263.64 64.18 263.64 64.18 273.45 10.63 273.45 10.63 206.24 2.34 206.24 2.34 206.12
         0.14 206.12 0.14 183.42 0.88 183.42 0.88 182.26 0.14 182.26 0.14 180.78 0.88 180.78 0.88 179.62 0.14 179.62 0.14 178.14
         0.88 178.14 0.88 176.98 0.14 176.98 0.14 175.5 0.88 175.5 0.88 174.34 0.14 174.34 0.14 0.14 149.86 0.14 ;
      LAYER M3 ;
      POLYGON 68.5 216.89 64.18 216.89 64.18 273.45 10.63 273.45 10.63 206.12 0.14 206.12 0.14 173.74 68.5 173.74 ;
      POLYGON 149.86 173.32 132.56 173.32 132.56 168.18 0.14 168.18 0.14 167.14 132.56 167.14 132.56 161.58 0.87 161.58 0.87 161.57 0.14 161.57 0.14 142.2
         0 142.2 0 141.6 0.14 141.6 0.14 136.92 0 136.92 0 136.32 0.14 136.32 0.14 111.84 0 111.84 0 111.24
         0.14 111.24 0.14 105.24 0 105.24 0 104.64 0.14 104.64 0.14 76.2 0 76.2 0 75.6 0.14 75.6 0.14 72.24
         0 72.24 0 71.64 0.14 71.64 0.14 45.84 0 45.84 0 45.24 0.14 45.24 0.14 41.88 0 41.88 0 41.28
         0.14 41.28 0.14 16.66 132.56 16.66 132.56 11.1 0.88 11.1 0.88 11.09 0.14 11.09 0.14 10.06 132.56 10.06 132.56 4.5
         0.88 4.5 0.88 4.49 0.14 4.49 0.14 0.14 149.86 0.14 ;
      LAYER M4 ;
      RECT 0.14 0.14 149.86 173.32 ;
      RECT 10.63 0.14 68.5 216.89 ;
      RECT 10.63 0.14 64.18 273.45 ;
      RECT 0.14 0.14 68.5 206.12 ;
  END
END pllclk

END LIBRARY
