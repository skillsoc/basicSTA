VERSION 5.4 ;
NAMESCASESENSITIVE ON ;

MACRO rom_512x16A
  CLASS RING ;
  FOREIGN rom_512x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 226.465 BY 184.645 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER M2 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER M3 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER M4 ;
      RECT 84.54 21.52 85.2 22.18 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER M2 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER M3 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER M4 ;
      RECT 80.44 21.52 81.1 22.18 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.039 ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER M2 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER M3 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER M4 ;
      RECT 76.34 21.52 77 22.18 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER M2 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER M3 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER M4 ;
      RECT 59.94 21.52 60.6 22.18 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER M2 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER M3 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER M4 ;
      RECT 55.84 21.52 56.5 22.18 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER M2 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER M3 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER M4 ;
      RECT 51.74 21.52 52.4 22.18 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER M2 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER M3 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER M4 ;
      RECT 43.54 21.52 44.2 22.18 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER M2 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER M3 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER M4 ;
      RECT 39.44 21.52 40.1 22.18 ;
      END
    END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER M2 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER M3 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER M4 ;
      RECT 35.34 21.52 36 22.18 ;
      END
    END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER M2 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER M3 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER M4 ;
      RECT 93.91 17.2 94.57 17.86 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER M1 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER M2 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER M3 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER M4 ;
      RECT 97.065 17.2 97.725 17.86 ;
      END
    END CLK
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER M2 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER M3 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER M4 ;
      RECT 118.055 17.2 118.715 17.86 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER M2 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER M3 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER M4 ;
      RECT 175.255 17.2 175.915 17.86 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER M2 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER M3 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER M4 ;
      RECT 180.375 17.2 181.035 17.86 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER M2 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER M3 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER M4 ;
      RECT 186.695 17.2 187.355 17.86 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER M2 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER M3 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER M4 ;
      RECT 191.815 17.2 192.475 17.86 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER M2 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER M3 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER M4 ;
      RECT 198.135 17.2 198.795 17.86 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER M2 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER M3 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER M4 ;
      RECT 203.255 17.2 203.915 17.86 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER M2 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER M3 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER M4 ;
      RECT 123.175 17.2 123.835 17.86 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER M2 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER M3 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER M4 ;
      RECT 129.495 17.2 130.155 17.86 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER M2 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER M3 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER M4 ;
      RECT 134.615 17.2 135.275 17.86 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER M2 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER M3 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER M4 ;
      RECT 140.935 17.2 141.595 17.86 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER M2 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER M3 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER M4 ;
      RECT 146.055 17.2 146.715 17.86 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER M2 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER M3 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER M4 ;
      RECT 152.375 17.2 153.035 17.86 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER M2 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER M3 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER M4 ;
      RECT 157.495 17.2 158.155 17.86 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER M2 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER M3 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER M4 ;
      RECT 163.815 17.2 164.475 17.86 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER M2 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER M3 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER M4 ;
      RECT 168.935 17.2 169.595 17.86 ;
      END
    END Q[9]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 226.465 176.645 0 184.645 ;
      LAYER M3 ;
      RECT 0 0 226.465 8 ;
      LAYER M4 ;
      RECT 218.465 0 226.465 184.645 ;
      LAYER M4 ;
      RECT 0 184.645 8 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 217.865 168.045 8.6 176.045 ;
      LAYER M3 ;
      RECT 8.6 8.6 217.865 16.6 ;
      LAYER M4 ;
      RECT 209.865 8.6 217.865 176.045 ;
      LAYER M4 ;
      RECT 8.6 176.045 16.6 8.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER V1 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER V2 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER V3 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER M1 ;
    POLYGON 17.2 167.445 17.2 21.52 35.16 21.52 35.16 22.36 36.18 22.36
      36.18 21.52 39.26 21.52 39.26 22.36 40.28 22.36 40.28 21.52 43.36 21.52
      43.36 22.36 44.38 22.36 44.38 21.52 51.56 21.52 51.56 22.36 52.58 22.36
      52.58 21.52 55.66 21.52 55.66 22.36 56.68 22.36 56.68 21.52 59.76 21.52
      59.76 22.36 60.78 22.36 60.78 21.52 76.16 21.52 76.16 22.36 77.18 22.36
      77.18 21.52 80.26 21.52 80.26 22.36 81.28 22.36 81.28 21.52 84.36 21.52
      84.36 22.36 85.38 22.36 85.38 21.52 91.99 21.52 91.99 17.2 93.73 17.2
      93.73 18.04 94.75 18.04 94.75 17.2 96.885 17.2 96.885 18.04
      97.905 18.04 97.905 17.2 117.875 17.2 117.875 18.04 118.895 18.04
      118.895 17.2 122.995 17.2 122.995 18.04 124.015 18.04 124.015 17.2
      129.315 17.2 129.315 18.04 130.335 18.04 130.335 17.2 134.435 17.2
      134.435 18.04 135.455 18.04 135.455 17.2 140.755 17.2 140.755 18.04
      141.775 18.04 141.775 17.2 145.875 17.2 145.875 18.04 146.895 18.04
      146.895 17.2 152.195 17.2 152.195 18.04 153.215 18.04 153.215 17.2
      157.315 17.2 157.315 18.04 158.335 18.04 158.335 17.2 163.635 17.2
      163.635 18.04 164.655 18.04 164.655 17.2 168.755 17.2 168.755 18.04
      169.775 18.04 169.775 17.2 175.075 17.2 175.075 18.04 176.095 18.04
      176.095 17.2 180.195 17.2 180.195 18.04 181.215 18.04 181.215 17.2
      186.515 17.2 186.515 18.04 187.535 18.04 187.535 17.2 191.635 17.2
      191.635 18.04 192.655 18.04 192.655 17.2 197.955 17.2 197.955 18.04
      198.975 18.04 198.975 17.2 203.075 17.2 203.075 18.04 204.095 18.04
      204.095 17.2 209.265 17.2 209.265 167.445 ;
    LAYER M2 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER M3 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER M4 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER M4 ;
    RECT 20.41 167.445 21.99 184.645 ;
    LAYER M4 ;
    RECT 24.57 167.445 26.15 184.645 ;
    LAYER M4 ;
    RECT 28.27 167.445 30.77 184.645 ;
    LAYER M4 ;
    RECT 36.47 167.445 38.97 184.645 ;
    LAYER M4 ;
    RECT 44.67 167.445 47.17 184.645 ;
    LAYER M4 ;
    RECT 52.87 167.445 55.37 184.645 ;
    LAYER M4 ;
    RECT 61.07 167.445 63.57 184.645 ;
    LAYER M4 ;
    RECT 69.27 167.445 71.77 184.645 ;
    LAYER M4 ;
    RECT 77.47 167.445 79.97 184.645 ;
    LAYER M4 ;
    RECT 85.67 167.445 88.17 184.645 ;
    LAYER M4 ;
    RECT 90.49 167.445 93.49 184.645 ;
    LAYER M4 ;
    RECT 97.63 167.445 100.63 184.645 ;
    LAYER M4 ;
    RECT 104.77 167.445 107.77 184.645 ;
    LAYER M4 ;
    RECT 110.85 167.445 112.65 184.645 ;
    LAYER M4 ;
    RECT 20.41 21.52 21.99 0 ;
    LAYER M4 ;
    RECT 24.57 21.52 26.15 0 ;
    LAYER M4 ;
    RECT 28.27 21.52 30.77 0 ;
    LAYER M4 ;
    RECT 36.47 21.52 38.97 0 ;
    LAYER M4 ;
    RECT 44.67 21.52 47.17 0 ;
    LAYER M4 ;
    RECT 52.87 21.52 55.37 0 ;
    LAYER M4 ;
    RECT 61.07 21.52 63.57 0 ;
    LAYER M4 ;
    RECT 69.27 21.52 71.77 0 ;
    LAYER M4 ;
    RECT 77.47 21.52 79.97 0 ;
    LAYER M4 ;
    RECT 85.67 21.52 88.17 0 ;
    LAYER M4 ;
    RECT 91.99 17.2 93.39 0 ;
    LAYER M4 ;
    RECT 98.415 17.2 99.815 0 ;
    LAYER M4 ;
    RECT 105 17.2 108 0 ;
    LAYER M4 ;
    RECT 110.85 17.2 112.65 0 ;
    LAYER M4 ;
    RECT 114.935 17.2 115.515 0 ;
    LAYER M4 ;
    RECT 117.015 17.2 117.595 0 ;
    LAYER M4 ;
    RECT 119.185 17.2 119.765 0 ;
    LAYER M4 ;
    RECT 122.125 17.2 122.705 0 ;
    LAYER M4 ;
    RECT 124.295 17.2 124.875 0 ;
    LAYER M4 ;
    RECT 126.375 17.2 126.955 0 ;
    LAYER M4 ;
    RECT 128.455 17.2 129.035 0 ;
    LAYER M4 ;
    RECT 130.625 17.2 131.205 0 ;
    LAYER M4 ;
    RECT 133.565 17.2 134.145 0 ;
    LAYER M4 ;
    RECT 135.735 17.2 136.315 0 ;
    LAYER M4 ;
    RECT 137.815 17.2 138.395 0 ;
    LAYER M4 ;
    RECT 139.895 17.2 140.475 0 ;
    LAYER M4 ;
    RECT 142.065 17.2 142.645 0 ;
    LAYER M4 ;
    RECT 145.005 17.2 145.585 0 ;
    LAYER M4 ;
    RECT 147.175 17.2 147.755 0 ;
    LAYER M4 ;
    RECT 149.255 17.2 149.835 0 ;
    LAYER M4 ;
    RECT 151.335 17.2 151.915 0 ;
    LAYER M4 ;
    RECT 153.505 17.2 154.085 0 ;
    LAYER M4 ;
    RECT 156.445 17.2 157.025 0 ;
    LAYER M4 ;
    RECT 158.615 17.2 159.195 0 ;
    LAYER M4 ;
    RECT 160.695 17.2 161.275 0 ;
    LAYER M4 ;
    RECT 162.775 17.2 163.355 0 ;
    LAYER M4 ;
    RECT 164.945 17.2 165.525 0 ;
    LAYER M4 ;
    RECT 167.885 17.2 168.465 0 ;
    LAYER M4 ;
    RECT 170.055 17.2 170.635 0 ;
    LAYER M4 ;
    RECT 172.135 17.2 172.715 0 ;
    LAYER M4 ;
    RECT 174.215 17.2 174.795 0 ;
    LAYER M4 ;
    RECT 176.385 17.2 176.965 0 ;
    LAYER M4 ;
    RECT 179.325 17.2 179.905 0 ;
    LAYER M4 ;
    RECT 181.495 17.2 182.075 0 ;
    LAYER M4 ;
    RECT 183.575 17.2 184.155 0 ;
    LAYER M4 ;
    RECT 185.655 17.2 186.235 0 ;
    LAYER M4 ;
    RECT 187.825 17.2 188.405 0 ;
    LAYER M4 ;
    RECT 190.765 17.2 191.345 0 ;
    LAYER M4 ;
    RECT 192.935 17.2 193.515 0 ;
    LAYER M4 ;
    RECT 195.015 17.2 195.595 0 ;
    LAYER M4 ;
    RECT 197.095 17.2 197.675 0 ;
    LAYER M4 ;
    RECT 199.265 17.2 199.845 0 ;
    LAYER M4 ;
    RECT 202.205 17.2 202.785 0 ;
    LAYER M4 ;
    RECT 204.375 17.2 204.955 0 ;
    LAYER M4 ;
    RECT 206.455 17.2 207.035 0 ;
    LAYER M3 ;
    RECT 209.265 21.085 226.465 22.485 ;
    LAYER M3 ;
    RECT 209.265 30.355 226.465 31.755 ;
    LAYER M3 ;
    RECT 209.265 32.615 226.465 34.015 ;
    LAYER M3 ;
    RECT 209.265 35.225 226.465 35.925 ;
    LAYER M3 ;
    RECT 209.265 40.26 226.465 42.74 ;
    LAYER M3 ;
    RECT 209.265 45.325 226.465 47.925 ;
    LAYER M3 ;
    RECT 209.265 50.515 226.465 51.755 ;
    LAYER M3 ;
    RECT 209.265 53.445 226.465 54.555 ;
    LAYER M3 ;
    RECT 209.265 57.13 226.465 57.83 ;
    LAYER M3 ;
    RECT 209.265 66.59 226.465 67.7 ;
    LAYER M3 ;
    RECT 209.265 72.31 226.465 74.11 ;
    LAYER M3 ;
    RECT 209.265 80.945 226.465 81.645 ;
    LAYER M3 ;
    RECT 209.265 84.125 226.465 85.925 ;
    LAYER M3 ;
    RECT 209.265 90.535 226.465 91.645 ;
    LAYER M3 ;
    RECT 209.265 100.045 226.465 100.745 ;
    LAYER M3 ;
    RECT 209.265 102.845 226.465 103.545 ;
    LAYER M3 ;
    RECT 209.265 109.675 226.465 112.075 ;
    LAYER M3 ;
    RECT 209.265 113.61 226.465 116.01 ;
    LAYER M3 ;
    RECT 17.2 24.88 0 25.58 ;
    LAYER M3 ;
    RECT 17.2 32.955 0 33.755 ;
    LAYER M3 ;
    RECT 17.2 35.055 0 35.755 ;
    LAYER M3 ;
    RECT 17.2 40.37 0 41.61 ;
    LAYER M3 ;
    RECT 17.2 43.96 0 46.56 ;
    LAYER M3 ;
    RECT 17.2 50.515 0 51.755 ;
    LAYER M3 ;
    RECT 17.2 53.445 0 54.555 ;
    LAYER M3 ;
    RECT 17.2 57.13 0 57.83 ;
    LAYER M3 ;
    RECT 17.2 66.59 0 67.7 ;
    LAYER M3 ;
    RECT 17.2 72.31 0 74.11 ;
    LAYER M3 ;
    RECT 17.2 80.885 0 81.585 ;
    LAYER M3 ;
    RECT 17.2 84.125 0 85.925 ;
    LAYER M3 ;
    RECT 17.2 90.535 0 91.645 ;
    LAYER M3 ;
    RECT 17.2 100.045 0 100.745 ;
    LAYER M3 ;
    RECT 17.2 109.675 0 112.075 ;
    LAYER M3 ;
    RECT 17.2 113.61 0 116.01 ;
    LAYER M3 ;
    RECT 17.2 124.62 0 125.32 ;
    LAYER M3 ;
    RECT 17.2 164.35 0 165.05 ;
    LAYER M4 ;
    RECT 22.49 167.445 24.07 176.045 ;
    LAYER M4 ;
    RECT 26.77 167.445 27.77 176.045 ;
    LAYER M4 ;
    RECT 32.37 167.445 34.87 176.045 ;
    LAYER M4 ;
    RECT 40.57 167.445 43.07 176.045 ;
    LAYER M4 ;
    RECT 48.77 167.445 51.27 176.045 ;
    LAYER M4 ;
    RECT 56.97 167.445 59.47 176.045 ;
    LAYER M4 ;
    RECT 65.17 167.445 67.67 176.045 ;
    LAYER M4 ;
    RECT 73.37 167.445 75.87 176.045 ;
    LAYER M4 ;
    RECT 81.57 167.445 84.07 176.045 ;
    LAYER M4 ;
    RECT 94.06 167.445 97.06 176.045 ;
    LAYER M4 ;
    RECT 101.2 167.445 104.2 176.045 ;
    LAYER M4 ;
    RECT 108.29 167.445 110.24 176.045 ;
    LAYER M4 ;
    RECT 113.67 167.445 115.07 176.045 ;
    LAYER M4 ;
    RECT 115.635 167.445 118.635 176.045 ;
    LAYER M4 ;
    RECT 119.755 167.445 121.755 176.045 ;
    LAYER M4 ;
    RECT 122.915 167.445 125.915 176.045 ;
    LAYER M4 ;
    RECT 127.075 167.445 130.075 176.045 ;
    LAYER M4 ;
    RECT 131.195 167.445 133.195 176.045 ;
    LAYER M4 ;
    RECT 134.355 167.445 137.355 176.045 ;
    LAYER M4 ;
    RECT 138.515 167.445 141.515 176.045 ;
    LAYER M4 ;
    RECT 142.635 167.445 144.635 176.045 ;
    LAYER M4 ;
    RECT 145.795 167.445 148.795 176.045 ;
    LAYER M4 ;
    RECT 149.955 167.445 152.955 176.045 ;
    LAYER M4 ;
    RECT 154.075 167.445 156.075 176.045 ;
    LAYER M4 ;
    RECT 157.235 167.445 160.235 176.045 ;
    LAYER M4 ;
    RECT 161.395 167.445 164.395 176.045 ;
    LAYER M4 ;
    RECT 165.515 167.445 167.515 176.045 ;
    LAYER M4 ;
    RECT 168.675 167.445 171.675 176.045 ;
    LAYER M4 ;
    RECT 172.835 167.445 175.835 176.045 ;
    LAYER M4 ;
    RECT 176.955 167.445 178.955 176.045 ;
    LAYER M4 ;
    RECT 180.115 167.445 183.115 176.045 ;
    LAYER M4 ;
    RECT 184.275 167.445 187.275 176.045 ;
    LAYER M4 ;
    RECT 188.395 167.445 190.395 176.045 ;
    LAYER M4 ;
    RECT 191.555 167.445 194.555 176.045 ;
    LAYER M4 ;
    RECT 195.715 167.445 198.715 176.045 ;
    LAYER M4 ;
    RECT 199.835 167.445 201.835 176.045 ;
    LAYER M4 ;
    RECT 202.995 167.445 205.995 176.045 ;
    LAYER M4 ;
    RECT 207.005 167.445 208.405 176.045 ;
    LAYER M4 ;
    RECT 22.49 21.52 24.07 8.6 ;
    LAYER M4 ;
    RECT 26.77 21.52 27.77 8.6 ;
    LAYER M4 ;
    RECT 32.37 21.52 34.87 8.6 ;
    LAYER M4 ;
    RECT 40.57 21.52 43.07 8.6 ;
    LAYER M4 ;
    RECT 48.77 21.52 51.27 8.6 ;
    LAYER M4 ;
    RECT 56.97 21.52 59.47 8.6 ;
    LAYER M4 ;
    RECT 65.17 21.52 67.67 8.6 ;
    LAYER M4 ;
    RECT 73.37 21.52 75.87 8.6 ;
    LAYER M4 ;
    RECT 81.57 21.52 84.07 8.6 ;
    LAYER M4 ;
    RECT 95.11 17.2 96.51 8.6 ;
    LAYER M4 ;
    RECT 101.54 17.2 104.54 8.6 ;
    LAYER M4 ;
    RECT 108.46 17.2 110.24 8.6 ;
    LAYER M4 ;
    RECT 113.205 17.2 114.405 8.6 ;
    LAYER M4 ;
    RECT 115.975 17.2 116.555 8.6 ;
    LAYER M4 ;
    RECT 120.345 17.2 121.545 8.6 ;
    LAYER M4 ;
    RECT 125.335 17.2 125.915 8.6 ;
    LAYER M4 ;
    RECT 127.415 17.2 127.995 8.6 ;
    LAYER M4 ;
    RECT 131.785 17.2 132.985 8.6 ;
    LAYER M4 ;
    RECT 136.775 17.2 137.355 8.6 ;
    LAYER M4 ;
    RECT 138.855 17.2 139.435 8.6 ;
    LAYER M4 ;
    RECT 143.225 17.2 144.425 8.6 ;
    LAYER M4 ;
    RECT 148.215 17.2 148.795 8.6 ;
    LAYER M4 ;
    RECT 150.295 17.2 150.875 8.6 ;
    LAYER M4 ;
    RECT 154.665 17.2 155.865 8.6 ;
    LAYER M4 ;
    RECT 159.655 17.2 160.235 8.6 ;
    LAYER M4 ;
    RECT 161.735 17.2 162.315 8.6 ;
    LAYER M4 ;
    RECT 166.105 17.2 167.305 8.6 ;
    LAYER M4 ;
    RECT 171.095 17.2 171.675 8.6 ;
    LAYER M4 ;
    RECT 173.175 17.2 173.755 8.6 ;
    LAYER M4 ;
    RECT 177.545 17.2 178.745 8.6 ;
    LAYER M4 ;
    RECT 182.535 17.2 183.115 8.6 ;
    LAYER M4 ;
    RECT 184.615 17.2 185.195 8.6 ;
    LAYER M4 ;
    RECT 188.985 17.2 190.185 8.6 ;
    LAYER M4 ;
    RECT 193.975 17.2 194.555 8.6 ;
    LAYER M4 ;
    RECT 196.055 17.2 196.635 8.6 ;
    LAYER M4 ;
    RECT 200.425 17.2 201.625 8.6 ;
    LAYER M4 ;
    RECT 205.415 17.2 205.995 8.6 ;
    LAYER M3 ;
    RECT 209.265 18.295 217.865 19.695 ;
    LAYER M3 ;
    RECT 209.265 23.685 217.865 25.085 ;
    LAYER M3 ;
    RECT 209.265 37.51 217.865 38.75 ;
    LAYER M3 ;
    RECT 209.265 48.825 217.865 49.625 ;
    LAYER M3 ;
    RECT 209.265 64.3 217.865 65.41 ;
    LAYER M3 ;
    RECT 209.265 68.16 217.865 68.86 ;
    LAYER M3 ;
    RECT 209.265 77.125 217.865 77.825 ;
    LAYER M3 ;
    RECT 209.265 82.105 217.865 83.215 ;
    LAYER M3 ;
    RECT 209.265 89.375 217.865 90.075 ;
    LAYER M3 ;
    RECT 209.265 92.765 217.865 93.875 ;
    LAYER M3 ;
    RECT 209.265 107.695 217.865 109.215 ;
    LAYER M3 ;
    RECT 209.265 118.19 217.865 120.19 ;
    LAYER M3 ;
    RECT 209.265 122.72 217.865 124.72 ;
    LAYER M3 ;
    RECT 209.265 125.22 217.865 127.22 ;
    LAYER M3 ;
    RECT 209.265 127.72 217.865 129.72 ;
    LAYER M3 ;
    RECT 209.265 130.22 217.865 132.22 ;
    LAYER M3 ;
    RECT 209.265 132.72 217.865 134.72 ;
    LAYER M3 ;
    RECT 209.265 135.22 217.865 137.22 ;
    LAYER M3 ;
    RECT 209.265 137.72 217.865 139.72 ;
    LAYER M3 ;
    RECT 209.265 140.22 217.865 142.22 ;
    LAYER M3 ;
    RECT 209.265 142.72 217.865 144.72 ;
    LAYER M3 ;
    RECT 209.265 145.22 217.865 147.22 ;
    LAYER M3 ;
    RECT 209.265 147.72 217.865 149.72 ;
    LAYER M3 ;
    RECT 209.265 150.22 217.865 152.22 ;
    LAYER M3 ;
    RECT 209.265 152.72 217.865 154.72 ;
    LAYER M3 ;
    RECT 209.265 155.22 217.865 157.22 ;
    LAYER M3 ;
    RECT 209.265 157.72 217.865 159.72 ;
    LAYER M3 ;
    RECT 209.265 160.22 217.865 162.22 ;
    LAYER M3 ;
    RECT 209.265 162.7 217.865 165.7 ;
    LAYER M3 ;
    RECT 17.2 27.815 8.6 28.615 ;
    LAYER M3 ;
    RECT 17.2 30.495 8.6 32.495 ;
    LAYER M3 ;
    RECT 17.2 36.215 8.6 37.455 ;
    LAYER M3 ;
    RECT 17.2 48.825 8.6 49.625 ;
    LAYER M3 ;
    RECT 17.2 64.3 8.6 65.41 ;
    LAYER M3 ;
    RECT 17.2 68.2 8.6 68.9 ;
    LAYER M3 ;
    RECT 17.2 77.125 8.6 77.825 ;
    LAYER M3 ;
    RECT 17.2 82.105 8.6 83.215 ;
    LAYER M3 ;
    RECT 17.2 89.335 8.6 90.035 ;
    LAYER M3 ;
    RECT 17.2 92.82 8.6 93.82 ;
    LAYER M3 ;
    RECT 17.2 107.815 8.6 109.215 ;
    LAYER M3 ;
    RECT 17.2 122.12 8.6 122.82 ;
    LAYER M3 ;
    RECT 17.2 127.12 8.6 127.82 ;
    LAYER M3 ;
    RECT 17.2 129.62 8.6 130.32 ;
    LAYER M3 ;
    RECT 17.2 132.12 8.6 132.82 ;
    LAYER M3 ;
    RECT 17.2 134.62 8.6 135.32 ;
    LAYER M3 ;
    RECT 17.2 137.12 8.6 137.82 ;
    LAYER M3 ;
    RECT 17.2 139.62 8.6 140.32 ;
    LAYER M3 ;
    RECT 17.2 142.12 8.6 142.82 ;
    LAYER M3 ;
    RECT 17.2 144.62 8.6 145.32 ;
    LAYER M3 ;
    RECT 17.2 147.12 8.6 147.82 ;
    LAYER M3 ;
    RECT 17.2 149.62 8.6 150.32 ;
    LAYER M3 ;
    RECT 17.2 152.12 8.6 152.82 ;
    LAYER M3 ;
    RECT 17.2 154.62 8.6 155.32 ;
    LAYER M3 ;
    RECT 17.2 157.12 8.6 157.82 ;
    LAYER M3 ;
    RECT 17.2 159.62 8.6 160.32 ;
    LAYER M3 ;
    RECT 17.2 162.12 8.6 162.82 ;
    END
  END rom_512x16A
END LIBRARY

