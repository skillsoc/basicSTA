VERSION 5.4 ;
NAMESCASESENSITIVE ON ;

MACRO ram_256x16A
  CLASS RING ;
  FOREIGN ram_256x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 256.485 BY 151.795 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 137.38 13.2 138.04 13.86 ;
      LAYER M2 ;
      RECT 137.38 13.2 138.04 13.86 ;
      LAYER M3 ;
      RECT 137.38 13.2 138.04 13.86 ;
      LAYER M4 ;
      RECT 137.38 13.2 138.04 13.86 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 131.26 13.2 131.92 13.86 ;
      LAYER M2 ;
      RECT 131.26 13.2 131.92 13.86 ;
      LAYER M3 ;
      RECT 131.26 13.2 131.92 13.86 ;
      LAYER M4 ;
      RECT 131.26 13.2 131.92 13.86 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 128.16 13.2 128.82 13.86 ;
      LAYER M2 ;
      RECT 128.16 13.2 128.82 13.86 ;
      LAYER M3 ;
      RECT 128.16 13.2 128.82 13.86 ;
      LAYER M4 ;
      RECT 128.16 13.2 128.82 13.86 ;
      END
    END A[2]
  PIN A[3]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 122.04 13.2 122.7 13.86 ;
      LAYER M2 ;
      RECT 122.04 13.2 122.7 13.86 ;
      LAYER M3 ;
      RECT 122.04 13.2 122.7 13.86 ;
      LAYER M4 ;
      RECT 122.04 13.2 122.7 13.86 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    ANTENNAGATEAREA  0.039 ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 119.02 13.2 119.68 13.86 ;
      LAYER M2 ;
      RECT 119.02 13.2 119.68 13.86 ;
      LAYER M3 ;
      RECT 119.02 13.2 119.68 13.86 ;
      LAYER M4 ;
      RECT 119.02 13.2 119.68 13.86 ;
      END
    END A[4]
  PIN A[5]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 115.92 13.2 116.58 13.86 ;
      LAYER M2 ;
      RECT 115.92 13.2 116.58 13.86 ;
      LAYER M3 ;
      RECT 115.92 13.2 116.58 13.86 ;
      LAYER M4 ;
      RECT 115.92 13.2 116.58 13.86 ;
      END
    END A[5]
  PIN A[6]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 109.8 13.2 110.46 13.86 ;
      LAYER M2 ;
      RECT 109.8 13.2 110.46 13.86 ;
      LAYER M3 ;
      RECT 109.8 13.2 110.46 13.86 ;
      LAYER M4 ;
      RECT 109.8 13.2 110.46 13.86 ;
      END
    END A[6]
  PIN A[7]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 106.78 13.2 107.44 13.86 ;
      LAYER M2 ;
      RECT 106.78 13.2 107.44 13.86 ;
      LAYER M3 ;
      RECT 106.78 13.2 107.44 13.86 ;
      LAYER M4 ;
      RECT 106.78 13.2 107.44 13.86 ;
      END
    END A[7]
  PIN CEN
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 143.195 13.2 143.855 13.86 ;
      LAYER M2 ;
      RECT 143.195 13.2 143.855 13.86 ;
      LAYER M3 ;
      RECT 143.195 13.2 143.855 13.86 ;
      LAYER M4 ;
      RECT 143.195 13.2 143.855 13.86 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    ANTENNAGATEAREA  0.039 ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
      RECT 152.94 13.2 153.6 13.86 ;
      LAYER M2 ;
      RECT 152.94 13.2 153.6 13.86 ;
      LAYER M3 ;
      RECT 152.94 13.2 153.6 13.86 ;
      LAYER M4 ;
      RECT 152.94 13.2 153.6 13.86 ;
      END
    END CLK
  PIN D[0]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 22.48 13.2 23.14 13.86 ;
      LAYER M2 ;
      RECT 22.48 13.2 23.14 13.86 ;
      LAYER M3 ;
      RECT 22.48 13.2 23.14 13.86 ;
      LAYER M4 ;
      RECT 22.48 13.2 23.14 13.86 ;
      END
    END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 181.685 13.2 182.345 13.86 ;
      LAYER M2 ;
      RECT 181.685 13.2 182.345 13.86 ;
      LAYER M3 ;
      RECT 181.685 13.2 182.345 13.86 ;
      LAYER M4 ;
      RECT 181.685 13.2 182.345 13.86 ;
      END
    END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 189.725 13.2 190.385 13.86 ;
      LAYER M2 ;
      RECT 189.725 13.2 190.385 13.86 ;
      LAYER M3 ;
      RECT 189.725 13.2 190.385 13.86 ;
      LAYER M4 ;
      RECT 189.725 13.2 190.385 13.86 ;
      END
    END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    ANTENNAGATEAREA  0.039 ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 204.025 13.2 204.685 13.86 ;
      LAYER M2 ;
      RECT 204.025 13.2 204.685 13.86 ;
      LAYER M3 ;
      RECT 204.025 13.2 204.685 13.86 ;
      LAYER M4 ;
      RECT 204.025 13.2 204.685 13.86 ;
      END
    END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 212.065 13.2 212.725 13.86 ;
      LAYER M2 ;
      RECT 212.065 13.2 212.725 13.86 ;
      LAYER M3 ;
      RECT 212.065 13.2 212.725 13.86 ;
      LAYER M4 ;
      RECT 212.065 13.2 212.725 13.86 ;
      END
    END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 225.305 13.2 225.965 13.86 ;
      LAYER M2 ;
      RECT 225.305 13.2 225.965 13.86 ;
      LAYER M3 ;
      RECT 225.305 13.2 225.965 13.86 ;
      LAYER M4 ;
      RECT 225.305 13.2 225.965 13.86 ;
      END
    END D[14]
  PIN D[15]
    ANTENNAGATEAREA  0.039 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 233.345 13.2 234.005 13.86 ;
      LAYER M2 ;
      RECT 233.345 13.2 234.005 13.86 ;
      LAYER M3 ;
      RECT 233.345 13.2 234.005 13.86 ;
      LAYER M4 ;
      RECT 233.345 13.2 234.005 13.86 ;
      END
    END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 30.52 13.2 31.18 13.86 ;
      LAYER M2 ;
      RECT 30.52 13.2 31.18 13.86 ;
      LAYER M3 ;
      RECT 30.52 13.2 31.18 13.86 ;
      LAYER M4 ;
      RECT 30.52 13.2 31.18 13.86 ;
      END
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 43.76 13.2 44.42 13.86 ;
      LAYER M2 ;
      RECT 43.76 13.2 44.42 13.86 ;
      LAYER M3 ;
      RECT 43.76 13.2 44.42 13.86 ;
      LAYER M4 ;
      RECT 43.76 13.2 44.42 13.86 ;
      END
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 51.8 13.2 52.46 13.86 ;
      LAYER M2 ;
      RECT 51.8 13.2 52.46 13.86 ;
      LAYER M3 ;
      RECT 51.8 13.2 52.46 13.86 ;
      LAYER M4 ;
      RECT 51.8 13.2 52.46 13.86 ;
      END
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 66.1 13.2 66.76 13.86 ;
      LAYER M2 ;
      RECT 66.1 13.2 66.76 13.86 ;
      LAYER M3 ;
      RECT 66.1 13.2 66.76 13.86 ;
      LAYER M4 ;
      RECT 66.1 13.2 66.76 13.86 ;
      END
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 74.14 13.2 74.8 13.86 ;
      LAYER M2 ;
      RECT 74.14 13.2 74.8 13.86 ;
      LAYER M3 ;
      RECT 74.14 13.2 74.8 13.86 ;
      LAYER M4 ;
      RECT 74.14 13.2 74.8 13.86 ;
      END
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 87.38 13.2 88.04 13.86 ;
      LAYER M2 ;
      RECT 87.38 13.2 88.04 13.86 ;
      LAYER M3 ;
      RECT 87.38 13.2 88.04 13.86 ;
      LAYER M4 ;
      RECT 87.38 13.2 88.04 13.86 ;
      END
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 95.42 13.2 96.08 13.86 ;
      LAYER M2 ;
      RECT 95.42 13.2 96.08 13.86 ;
      LAYER M3 ;
      RECT 95.42 13.2 96.08 13.86 ;
      LAYER M4 ;
      RECT 95.42 13.2 96.08 13.86 ;
      END
    END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 160.405 13.2 161.065 13.86 ;
      LAYER M2 ;
      RECT 160.405 13.2 161.065 13.86 ;
      LAYER M3 ;
      RECT 160.405 13.2 161.065 13.86 ;
      LAYER M4 ;
      RECT 160.405 13.2 161.065 13.86 ;
      END
    END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA  0.039 ;
    PORT
      LAYER M1 ;
      RECT 168.445 13.2 169.105 13.86 ;
      LAYER M2 ;
      RECT 168.445 13.2 169.105 13.86 ;
      LAYER M3 ;
      RECT 168.445 13.2 169.105 13.86 ;
      LAYER M4 ;
      RECT 168.445 13.2 169.105 13.86 ;
      END
    END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 25.06 13.2 25.72 13.86 ;
      LAYER M2 ;
      RECT 25.06 13.2 25.72 13.86 ;
      LAYER M3 ;
      RECT 25.06 13.2 25.72 13.86 ;
      LAYER M4 ;
      RECT 25.06 13.2 25.72 13.86 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 184.265 13.2 184.925 13.86 ;
      LAYER M2 ;
      RECT 184.265 13.2 184.925 13.86 ;
      LAYER M3 ;
      RECT 184.265 13.2 184.925 13.86 ;
      LAYER M4 ;
      RECT 184.265 13.2 184.925 13.86 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 187.145 13.2 187.805 13.86 ;
      LAYER M2 ;
      RECT 187.145 13.2 187.805 13.86 ;
      LAYER M3 ;
      RECT 187.145 13.2 187.805 13.86 ;
      LAYER M4 ;
      RECT 187.145 13.2 187.805 13.86 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 206.605 13.2 207.265 13.86 ;
      LAYER M2 ;
      RECT 206.605 13.2 207.265 13.86 ;
      LAYER M3 ;
      RECT 206.605 13.2 207.265 13.86 ;
      LAYER M4 ;
      RECT 206.605 13.2 207.265 13.86 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 209.485 13.2 210.145 13.86 ;
      LAYER M2 ;
      RECT 209.485 13.2 210.145 13.86 ;
      LAYER M3 ;
      RECT 209.485 13.2 210.145 13.86 ;
      LAYER M4 ;
      RECT 209.485 13.2 210.145 13.86 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 227.885 13.2 228.545 13.86 ;
      LAYER M2 ;
      RECT 227.885 13.2 228.545 13.86 ;
      LAYER M3 ;
      RECT 227.885 13.2 228.545 13.86 ;
      LAYER M4 ;
      RECT 227.885 13.2 228.545 13.86 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 230.765 13.2 231.425 13.86 ;
      LAYER M2 ;
      RECT 230.765 13.2 231.425 13.86 ;
      LAYER M3 ;
      RECT 230.765 13.2 231.425 13.86 ;
      LAYER M4 ;
      RECT 230.765 13.2 231.425 13.86 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 27.94 13.2 28.6 13.86 ;
      LAYER M2 ;
      RECT 27.94 13.2 28.6 13.86 ;
      LAYER M3 ;
      RECT 27.94 13.2 28.6 13.86 ;
      LAYER M4 ;
      RECT 27.94 13.2 28.6 13.86 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 46.34 13.2 47 13.86 ;
      LAYER M2 ;
      RECT 46.34 13.2 47 13.86 ;
      LAYER M3 ;
      RECT 46.34 13.2 47 13.86 ;
      LAYER M4 ;
      RECT 46.34 13.2 47 13.86 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 49.22 13.2 49.88 13.86 ;
      LAYER M2 ;
      RECT 49.22 13.2 49.88 13.86 ;
      LAYER M3 ;
      RECT 49.22 13.2 49.88 13.86 ;
      LAYER M4 ;
      RECT 49.22 13.2 49.88 13.86 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 68.68 13.2 69.34 13.86 ;
      LAYER M2 ;
      RECT 68.68 13.2 69.34 13.86 ;
      LAYER M3 ;
      RECT 68.68 13.2 69.34 13.86 ;
      LAYER M4 ;
      RECT 68.68 13.2 69.34 13.86 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 71.56 13.2 72.22 13.86 ;
      LAYER M2 ;
      RECT 71.56 13.2 72.22 13.86 ;
      LAYER M3 ;
      RECT 71.56 13.2 72.22 13.86 ;
      LAYER M4 ;
      RECT 71.56 13.2 72.22 13.86 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 89.96 13.2 90.62 13.86 ;
      LAYER M2 ;
      RECT 89.96 13.2 90.62 13.86 ;
      LAYER M3 ;
      RECT 89.96 13.2 90.62 13.86 ;
      LAYER M4 ;
      RECT 89.96 13.2 90.62 13.86 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 92.84 13.2 93.5 13.86 ;
      LAYER M2 ;
      RECT 92.84 13.2 93.5 13.86 ;
      LAYER M3 ;
      RECT 92.84 13.2 93.5 13.86 ;
      LAYER M4 ;
      RECT 92.84 13.2 93.5 13.86 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 162.985 13.2 163.645 13.86 ;
      LAYER M2 ;
      RECT 162.985 13.2 163.645 13.86 ;
      LAYER M3 ;
      RECT 162.985 13.2 163.645 13.86 ;
      LAYER M4 ;
      RECT 162.985 13.2 163.645 13.86 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 165.865 13.2 166.525 13.86 ;
      LAYER M2 ;
      RECT 165.865 13.2 166.525 13.86 ;
      LAYER M3 ;
      RECT 165.865 13.2 166.525 13.86 ;
      LAYER M4 ;
      RECT 165.865 13.2 166.525 13.86 ;
      END
    END Q[9]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 149.24 13.2 149.9 13.86 ;
      LAYER M2 ;
      RECT 149.24 13.2 149.9 13.86 ;
      LAYER M3 ;
      RECT 149.24 13.2 149.9 13.86 ;
      LAYER M4 ;
      RECT 149.24 13.2 149.9 13.86 ;
      END
    END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 256.485 145.795 0 151.795 ;
      LAYER M3 ;
      RECT 0 0 256.485 6 ;
      LAYER M4 ;
      RECT 250.485 0 256.485 151.795 ;
      LAYER M4 ;
      RECT 0 151.795 6 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 249.885 139.195 6.6 145.195 ;
      LAYER M3 ;
      RECT 6.6 6.6 249.885 12.6 ;
      LAYER M4 ;
      RECT 243.885 6.6 249.885 145.195 ;
      LAYER M4 ;
      RECT 6.6 145.195 12.6 6.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 13.2 13.2 243.285 138.595 ;
    LAYER V1 ;
    RECT 13.2 13.2 243.285 138.595 ;
    LAYER V2 ;
    RECT 13.2 13.2 243.285 138.595 ;
    LAYER V3 ;
    RECT 13.2 13.2 243.285 138.595 ;
    LAYER M1 ;
    POLYGON 13.2 138.595 13.2 13.2 22.3 13.2 22.3 14.04 23.32 14.04
      23.32 13.2 24.88 13.2 24.88 14.04 25.9 14.04 25.9 13.2 27.76 13.2
      27.76 14.04 28.78 14.04 28.78 13.2 30.34 13.2 30.34 14.04 31.36 14.04
      31.36 13.2 43.58 13.2 43.58 14.04 44.6 14.04 44.6 13.2 46.16 13.2
      46.16 14.04 47.18 14.04 47.18 13.2 49.04 13.2 49.04 14.04 50.06 14.04
      50.06 13.2 51.62 13.2 51.62 14.04 52.64 14.04 52.64 13.2 65.92 13.2
      65.92 14.04 66.94 14.04 66.94 13.2 68.5 13.2 68.5 14.04 69.52 14.04
      69.52 13.2 71.38 13.2 71.38 14.04 72.4 14.04 72.4 13.2 73.96 13.2
      73.96 14.04 74.98 14.04 74.98 13.2 87.2 13.2 87.2 14.04 88.22 14.04
      88.22 13.2 89.78 13.2 89.78 14.04 90.8 14.04 90.8 13.2 92.66 13.2
      92.66 14.04 93.68 14.04 93.68 13.2 95.24 13.2 95.24 14.04 96.26 14.04
      96.26 13.2 106.6 13.2 106.6 14.04 107.62 14.04 107.62 13.2 109.62 13.2
      109.62 14.04 110.64 14.04 110.64 13.2 115.74 13.2 115.74 14.04
      116.76 14.04 116.76 13.2 118.84 13.2 118.84 14.04 119.86 14.04
      119.86 13.2 121.86 13.2 121.86 14.04 122.88 14.04 122.88 13.2
      127.98 13.2 127.98 14.04 129 14.04 129 13.2 131.08 13.2 131.08 14.04
      132.1 14.04 132.1 13.2 137.2 13.2 137.2 14.04 138.22 14.04 138.22 13.2
      143.015 13.2 143.015 14.04 144.035 14.04 144.035 13.2 149.06 13.2
      149.06 14.04 150.08 14.04 150.08 13.2 152.76 13.2 152.76 14.04
      153.78 14.04 153.78 13.2 160.225 13.2 160.225 14.04 161.245 14.04
      161.245 13.2 162.805 13.2 162.805 14.04 163.825 14.04 163.825 13.2
      165.685 13.2 165.685 14.04 166.705 14.04 166.705 13.2 168.265 13.2
      168.265 14.04 169.285 14.04 169.285 13.2 181.505 13.2 181.505 14.04
      182.525 14.04 182.525 13.2 184.085 13.2 184.085 14.04 185.105 14.04
      185.105 13.2 186.965 13.2 186.965 14.04 187.985 14.04 187.985 13.2
      189.545 13.2 189.545 14.04 190.565 14.04 190.565 13.2 203.845 13.2
      203.845 14.04 204.865 14.04 204.865 13.2 206.425 13.2 206.425 14.04
      207.445 14.04 207.445 13.2 209.305 13.2 209.305 14.04 210.325 14.04
      210.325 13.2 211.885 13.2 211.885 14.04 212.905 14.04 212.905 13.2
      225.125 13.2 225.125 14.04 226.145 14.04 226.145 13.2 227.705 13.2
      227.705 14.04 228.725 14.04 228.725 13.2 230.585 13.2 230.585 14.04
      231.605 14.04 231.605 13.2 233.165 13.2 233.165 14.04 234.185 14.04
      234.185 13.2 243.285 13.2 243.285 138.595 ;
    LAYER M2 ;
    POLYGON 13.2 138.595 13.2 13.2 22.27 13.2 22.27 14.07 23.35 14.07
      23.35 13.2 24.85 13.2 24.85 14.07 25.93 14.07 25.93 13.2 27.73 13.2
      27.73 14.07 28.81 14.07 28.81 13.2 30.31 13.2 30.31 14.07 31.39 14.07
      31.39 13.2 43.55 13.2 43.55 14.07 44.63 14.07 44.63 13.2 46.13 13.2
      46.13 14.07 47.21 14.07 47.21 13.2 49.01 13.2 49.01 14.07 50.09 14.07
      50.09 13.2 51.59 13.2 51.59 14.07 52.67 14.07 52.67 13.2 65.89 13.2
      65.89 14.07 66.97 14.07 66.97 13.2 68.47 13.2 68.47 14.07 69.55 14.07
      69.55 13.2 71.35 13.2 71.35 14.07 72.43 14.07 72.43 13.2 73.93 13.2
      73.93 14.07 75.01 14.07 75.01 13.2 87.17 13.2 87.17 14.07 88.25 14.07
      88.25 13.2 89.75 13.2 89.75 14.07 90.83 14.07 90.83 13.2 92.63 13.2
      92.63 14.07 93.71 14.07 93.71 13.2 95.21 13.2 95.21 14.07 96.29 14.07
      96.29 13.2 106.57 13.2 106.57 14.07 107.65 14.07 107.65 13.2
      109.59 13.2 109.59 14.07 110.67 14.07 110.67 13.2 115.71 13.2
      115.71 14.07 116.79 14.07 116.79 13.2 118.81 13.2 118.81 14.07
      119.89 14.07 119.89 13.2 121.83 13.2 121.83 14.07 122.91 14.07
      122.91 13.2 127.95 13.2 127.95 14.07 129.03 14.07 129.03 13.2
      131.05 13.2 131.05 14.07 132.13 14.07 132.13 13.2 137.17 13.2
      137.17 14.07 138.25 14.07 138.25 13.2 142.985 13.2 142.985 14.07
      144.065 14.07 144.065 13.2 149.03 13.2 149.03 14.07 150.11 14.07
      150.11 13.2 152.73 13.2 152.73 14.07 153.81 14.07 153.81 13.2
      160.195 13.2 160.195 14.07 161.275 14.07 161.275 13.2 162.775 13.2
      162.775 14.07 163.855 14.07 163.855 13.2 165.655 13.2 165.655 14.07
      166.735 14.07 166.735 13.2 168.235 13.2 168.235 14.07 169.315 14.07
      169.315 13.2 181.475 13.2 181.475 14.07 182.555 14.07 182.555 13.2
      184.055 13.2 184.055 14.07 185.135 14.07 185.135 13.2 186.935 13.2
      186.935 14.07 188.015 14.07 188.015 13.2 189.515 13.2 189.515 14.07
      190.595 14.07 190.595 13.2 203.815 13.2 203.815 14.07 204.895 14.07
      204.895 13.2 206.395 13.2 206.395 14.07 207.475 14.07 207.475 13.2
      209.275 13.2 209.275 14.07 210.355 14.07 210.355 13.2 211.855 13.2
      211.855 14.07 212.935 14.07 212.935 13.2 225.095 13.2 225.095 14.07
      226.175 14.07 226.175 13.2 227.675 13.2 227.675 14.07 228.755 14.07
      228.755 13.2 230.555 13.2 230.555 14.07 231.635 14.07 231.635 13.2
      233.135 13.2 233.135 14.07 234.215 14.07 234.215 13.2 243.285 13.2
      243.285 138.595 ;
    LAYER M3 ;
    POLYGON 13.2 138.595 13.2 13.2 22.27 13.2 22.27 14.07 23.35 14.07
      23.35 13.2 24.85 13.2 24.85 14.07 25.93 14.07 25.93 13.2 27.73 13.2
      27.73 14.07 28.81 14.07 28.81 13.2 30.31 13.2 30.31 14.07 31.39 14.07
      31.39 13.2 43.55 13.2 43.55 14.07 44.63 14.07 44.63 13.2 46.13 13.2
      46.13 14.07 47.21 14.07 47.21 13.2 49.01 13.2 49.01 14.07 50.09 14.07
      50.09 13.2 51.59 13.2 51.59 14.07 52.67 14.07 52.67 13.2 65.89 13.2
      65.89 14.07 66.97 14.07 66.97 13.2 68.47 13.2 68.47 14.07 69.55 14.07
      69.55 13.2 71.35 13.2 71.35 14.07 72.43 14.07 72.43 13.2 73.93 13.2
      73.93 14.07 75.01 14.07 75.01 13.2 87.17 13.2 87.17 14.07 88.25 14.07
      88.25 13.2 89.75 13.2 89.75 14.07 90.83 14.07 90.83 13.2 92.63 13.2
      92.63 14.07 93.71 14.07 93.71 13.2 95.21 13.2 95.21 14.07 96.29 14.07
      96.29 13.2 106.57 13.2 106.57 14.07 107.65 14.07 107.65 13.2
      109.59 13.2 109.59 14.07 110.67 14.07 110.67 13.2 115.71 13.2
      115.71 14.07 116.79 14.07 116.79 13.2 118.81 13.2 118.81 14.07
      119.89 14.07 119.89 13.2 121.83 13.2 121.83 14.07 122.91 14.07
      122.91 13.2 127.95 13.2 127.95 14.07 129.03 14.07 129.03 13.2
      131.05 13.2 131.05 14.07 132.13 14.07 132.13 13.2 137.17 13.2
      137.17 14.07 138.25 14.07 138.25 13.2 142.985 13.2 142.985 14.07
      144.065 14.07 144.065 13.2 149.03 13.2 149.03 14.07 150.11 14.07
      150.11 13.2 152.73 13.2 152.73 14.07 153.81 14.07 153.81 13.2
      160.195 13.2 160.195 14.07 161.275 14.07 161.275 13.2 162.775 13.2
      162.775 14.07 163.855 14.07 163.855 13.2 165.655 13.2 165.655 14.07
      166.735 14.07 166.735 13.2 168.235 13.2 168.235 14.07 169.315 14.07
      169.315 13.2 181.475 13.2 181.475 14.07 182.555 14.07 182.555 13.2
      184.055 13.2 184.055 14.07 185.135 14.07 185.135 13.2 186.935 13.2
      186.935 14.07 188.015 14.07 188.015 13.2 189.515 13.2 189.515 14.07
      190.595 14.07 190.595 13.2 203.815 13.2 203.815 14.07 204.895 14.07
      204.895 13.2 206.395 13.2 206.395 14.07 207.475 14.07 207.475 13.2
      209.275 13.2 209.275 14.07 210.355 14.07 210.355 13.2 211.855 13.2
      211.855 14.07 212.935 14.07 212.935 13.2 225.095 13.2 225.095 14.07
      226.175 14.07 226.175 13.2 227.675 13.2 227.675 14.07 228.755 14.07
      228.755 13.2 230.555 13.2 230.555 14.07 231.635 14.07 231.635 13.2
      233.135 13.2 233.135 14.07 234.215 14.07 234.215 13.2 243.285 13.2
      243.285 138.595 ;
    LAYER M4 ;
    POLYGON 13.2 138.595 13.2 13.2 22.27 13.2 22.27 14.07 23.35 14.07
      23.35 13.2 24.85 13.2 24.85 14.07 25.93 14.07 25.93 13.2 27.73 13.2
      27.73 14.07 28.81 14.07 28.81 13.2 30.31 13.2 30.31 14.07 31.39 14.07
      31.39 13.2 43.55 13.2 43.55 14.07 44.63 14.07 44.63 13.2 46.13 13.2
      46.13 14.07 47.21 14.07 47.21 13.2 49.01 13.2 49.01 14.07 50.09 14.07
      50.09 13.2 51.59 13.2 51.59 14.07 52.67 14.07 52.67 13.2 65.89 13.2
      65.89 14.07 66.97 14.07 66.97 13.2 68.47 13.2 68.47 14.07 69.55 14.07
      69.55 13.2 71.35 13.2 71.35 14.07 72.43 14.07 72.43 13.2 73.93 13.2
      73.93 14.07 75.01 14.07 75.01 13.2 87.17 13.2 87.17 14.07 88.25 14.07
      88.25 13.2 89.75 13.2 89.75 14.07 90.83 14.07 90.83 13.2 92.63 13.2
      92.63 14.07 93.71 14.07 93.71 13.2 95.21 13.2 95.21 14.07 96.29 14.07
      96.29 13.2 106.57 13.2 106.57 14.07 107.65 14.07 107.65 13.2
      109.59 13.2 109.59 14.07 110.67 14.07 110.67 13.2 115.71 13.2
      115.71 14.07 116.79 14.07 116.79 13.2 118.81 13.2 118.81 14.07
      119.89 14.07 119.89 13.2 121.83 13.2 121.83 14.07 122.91 14.07
      122.91 13.2 127.95 13.2 127.95 14.07 129.03 14.07 129.03 13.2
      131.05 13.2 131.05 14.07 132.13 14.07 132.13 13.2 137.17 13.2
      137.17 14.07 138.25 14.07 138.25 13.2 142.985 13.2 142.985 14.07
      144.065 14.07 144.065 13.2 149.03 13.2 149.03 14.07 150.11 14.07
      150.11 13.2 152.73 13.2 152.73 14.07 153.81 14.07 153.81 13.2
      160.195 13.2 160.195 14.07 161.275 14.07 161.275 13.2 162.775 13.2
      162.775 14.07 163.855 14.07 163.855 13.2 165.655 13.2 165.655 14.07
      166.735 14.07 166.735 13.2 168.235 13.2 168.235 14.07 169.315 14.07
      169.315 13.2 181.475 13.2 181.475 14.07 182.555 14.07 182.555 13.2
      184.055 13.2 184.055 14.07 185.135 14.07 185.135 13.2 186.935 13.2
      186.935 14.07 188.015 14.07 188.015 13.2 189.515 13.2 189.515 14.07
      190.595 14.07 190.595 13.2 203.815 13.2 203.815 14.07 204.895 14.07
      204.895 13.2 206.395 13.2 206.395 14.07 207.475 14.07 207.475 13.2
      209.275 13.2 209.275 14.07 210.355 14.07 210.355 13.2 211.855 13.2
      211.855 14.07 212.935 14.07 212.935 13.2 225.095 13.2 225.095 14.07
      226.175 14.07 226.175 13.2 227.675 13.2 227.675 14.07 228.755 14.07
      228.755 13.2 230.555 13.2 230.555 14.07 231.635 14.07 231.635 13.2
      233.135 13.2 233.135 14.07 234.215 14.07 234.215 13.2 243.285 13.2
      243.285 138.595 ;
    LAYER M4 ;
    RECT 17.775 138.595 18.595 151.795 ;
    LAYER M4 ;
    RECT 19.105 138.595 19.925 151.795 ;
    LAYER M4 ;
    RECT 23.095 138.595 23.915 151.795 ;
    LAYER M4 ;
    RECT 24.425 138.595 25.245 151.795 ;
    LAYER M4 ;
    RECT 28.415 138.595 29.235 151.795 ;
    LAYER M4 ;
    RECT 29.745 138.595 30.565 151.795 ;
    LAYER M4 ;
    RECT 33.735 138.595 34.555 151.795 ;
    LAYER M4 ;
    RECT 35.065 138.595 35.885 151.795 ;
    LAYER M4 ;
    RECT 39.055 138.595 39.875 151.795 ;
    LAYER M4 ;
    RECT 40.385 138.595 41.205 151.795 ;
    LAYER M4 ;
    RECT 44.375 138.595 45.195 151.795 ;
    LAYER M4 ;
    RECT 45.705 138.595 46.525 151.795 ;
    LAYER M4 ;
    RECT 49.695 138.595 50.515 151.795 ;
    LAYER M4 ;
    RECT 51.025 138.595 51.845 151.795 ;
    LAYER M4 ;
    RECT 55.015 138.595 55.835 151.795 ;
    LAYER M4 ;
    RECT 56.345 138.595 57.165 151.795 ;
    LAYER M4 ;
    RECT 61.395 138.595 62.215 151.795 ;
    LAYER M4 ;
    RECT 62.725 138.595 63.545 151.795 ;
    LAYER M4 ;
    RECT 66.715 138.595 67.535 151.795 ;
    LAYER M4 ;
    RECT 68.045 138.595 68.865 151.795 ;
    LAYER M4 ;
    RECT 72.035 138.595 72.855 151.795 ;
    LAYER M4 ;
    RECT 73.365 138.595 74.185 151.795 ;
    LAYER M4 ;
    RECT 77.355 138.595 78.175 151.795 ;
    LAYER M4 ;
    RECT 78.685 138.595 79.505 151.795 ;
    LAYER M4 ;
    RECT 82.675 138.595 83.495 151.795 ;
    LAYER M4 ;
    RECT 84.005 138.595 84.825 151.795 ;
    LAYER M4 ;
    RECT 87.995 138.595 88.815 151.795 ;
    LAYER M4 ;
    RECT 89.325 138.595 90.145 151.795 ;
    LAYER M4 ;
    RECT 93.315 138.595 94.135 151.795 ;
    LAYER M4 ;
    RECT 94.645 138.595 95.465 151.795 ;
    LAYER M4 ;
    RECT 98.635 138.595 99.455 151.795 ;
    LAYER M4 ;
    RECT 99.965 138.595 100.785 151.795 ;
    LAYER M4 ;
    RECT 103.715 138.595 104.975 151.795 ;
    LAYER M4 ;
    RECT 105.79 138.595 106.85 151.795 ;
    LAYER M4 ;
    RECT 108.85 138.595 109.91 151.795 ;
    LAYER M4 ;
    RECT 111.91 138.595 112.97 151.795 ;
    LAYER M4 ;
    RECT 114.97 138.595 116.03 151.795 ;
    LAYER M4 ;
    RECT 118.03 138.595 119.09 151.795 ;
    LAYER M4 ;
    RECT 121.09 138.595 122.15 151.795 ;
    LAYER M4 ;
    RECT 124.15 138.595 125.21 151.795 ;
    LAYER M4 ;
    RECT 127.21 138.595 128.27 151.795 ;
    LAYER M4 ;
    RECT 130.27 138.595 131.33 151.795 ;
    LAYER M4 ;
    RECT 133.33 138.595 134.39 151.795 ;
    LAYER M4 ;
    RECT 136.39 138.595 137.45 151.795 ;
    LAYER M4 ;
    RECT 139.835 138.595 141.095 151.795 ;
    LAYER M4 ;
    RECT 143.915 138.595 145.175 151.795 ;
    LAYER M4 ;
    RECT 147.995 138.595 149.255 151.795 ;
    LAYER M4 ;
    RECT 151.98 138.595 152.8 151.795 ;
    LAYER M4 ;
    RECT 155.7 138.595 156.52 151.795 ;
    LAYER M4 ;
    RECT 157.03 138.595 157.85 151.795 ;
    LAYER M4 ;
    RECT 161.02 138.595 161.84 151.795 ;
    LAYER M4 ;
    RECT 162.35 138.595 163.17 151.795 ;
    LAYER M4 ;
    RECT 166.34 138.595 167.16 151.795 ;
    LAYER M4 ;
    RECT 167.67 138.595 168.49 151.795 ;
    LAYER M4 ;
    RECT 171.66 138.595 172.48 151.795 ;
    LAYER M4 ;
    RECT 172.99 138.595 173.81 151.795 ;
    LAYER M4 ;
    RECT 176.98 138.595 177.8 151.795 ;
    LAYER M4 ;
    RECT 178.31 138.595 179.13 151.795 ;
    LAYER M4 ;
    RECT 182.3 138.595 183.12 151.795 ;
    LAYER M4 ;
    RECT 183.63 138.595 184.45 151.795 ;
    LAYER M4 ;
    RECT 187.62 138.595 188.44 151.795 ;
    LAYER M4 ;
    RECT 188.95 138.595 189.77 151.795 ;
    LAYER M4 ;
    RECT 192.94 138.595 193.76 151.795 ;
    LAYER M4 ;
    RECT 194.27 138.595 195.09 151.795 ;
    LAYER M4 ;
    RECT 199.32 138.595 200.14 151.795 ;
    LAYER M4 ;
    RECT 200.65 138.595 201.47 151.795 ;
    LAYER M4 ;
    RECT 204.64 138.595 205.46 151.795 ;
    LAYER M4 ;
    RECT 205.97 138.595 206.79 151.795 ;
    LAYER M4 ;
    RECT 209.96 138.595 210.78 151.795 ;
    LAYER M4 ;
    RECT 211.29 138.595 212.11 151.795 ;
    LAYER M4 ;
    RECT 215.28 138.595 216.1 151.795 ;
    LAYER M4 ;
    RECT 216.61 138.595 217.43 151.795 ;
    LAYER M4 ;
    RECT 220.6 138.595 221.42 151.795 ;
    LAYER M4 ;
    RECT 221.93 138.595 222.75 151.795 ;
    LAYER M4 ;
    RECT 225.92 138.595 226.74 151.795 ;
    LAYER M4 ;
    RECT 227.25 138.595 228.07 151.795 ;
    LAYER M4 ;
    RECT 231.24 138.595 232.06 151.795 ;
    LAYER M4 ;
    RECT 232.57 138.595 233.39 151.795 ;
    LAYER M4 ;
    RECT 236.56 138.595 237.38 151.795 ;
    LAYER M4 ;
    RECT 237.89 138.595 238.71 151.795 ;
    LAYER M4 ;
    RECT 18.96 13.2 20.26 0 ;
    LAYER M4 ;
    RECT 23.6 13.2 24.6 0 ;
    LAYER M4 ;
    RECT 29.06 13.2 30.06 0 ;
    LAYER M4 ;
    RECT 33.4 13.2 34.7 0 ;
    LAYER M4 ;
    RECT 40.24 13.2 41.54 0 ;
    LAYER M4 ;
    RECT 44.88 13.2 45.88 0 ;
    LAYER M4 ;
    RECT 50.34 13.2 51.34 0 ;
    LAYER M4 ;
    RECT 54.68 13.2 55.98 0 ;
    LAYER M4 ;
    RECT 62.58 13.2 63.88 0 ;
    LAYER M4 ;
    RECT 67.22 13.2 68.22 0 ;
    LAYER M4 ;
    RECT 72.68 13.2 73.68 0 ;
    LAYER M4 ;
    RECT 77.02 13.2 78.32 0 ;
    LAYER M4 ;
    RECT 83.86 13.2 85.16 0 ;
    LAYER M4 ;
    RECT 88.5 13.2 89.5 0 ;
    LAYER M4 ;
    RECT 93.96 13.2 94.96 0 ;
    LAYER M4 ;
    RECT 98.3 13.2 99.6 0 ;
    LAYER M4 ;
    RECT 103.175 13.2 104.435 0 ;
    LAYER M4 ;
    RECT 107.99 13.2 109.25 0 ;
    LAYER M4 ;
    RECT 114.11 13.2 115.37 0 ;
    LAYER M4 ;
    RECT 120.23 13.2 121.49 0 ;
    LAYER M4 ;
    RECT 126.35 13.2 127.61 0 ;
    LAYER M4 ;
    RECT 132.47 13.2 133.73 0 ;
    LAYER M4 ;
    RECT 138.59 13.2 139.85 0 ;
    LAYER M4 ;
    RECT 140.31 13.2 141.01 0 ;
    LAYER M4 ;
    RECT 144.315 13.2 145.135 0 ;
    LAYER M4 ;
    RECT 147.78 13.2 148.78 0 ;
    LAYER M4 ;
    RECT 156.885 13.2 158.185 0 ;
    LAYER M4 ;
    RECT 161.525 13.2 162.525 0 ;
    LAYER M4 ;
    RECT 166.985 13.2 167.985 0 ;
    LAYER M4 ;
    RECT 171.325 13.2 172.625 0 ;
    LAYER M4 ;
    RECT 178.165 13.2 179.465 0 ;
    LAYER M4 ;
    RECT 182.805 13.2 183.805 0 ;
    LAYER M4 ;
    RECT 188.265 13.2 189.265 0 ;
    LAYER M4 ;
    RECT 192.605 13.2 193.905 0 ;
    LAYER M4 ;
    RECT 200.505 13.2 201.805 0 ;
    LAYER M4 ;
    RECT 205.145 13.2 206.145 0 ;
    LAYER M4 ;
    RECT 210.605 13.2 211.605 0 ;
    LAYER M4 ;
    RECT 214.945 13.2 216.245 0 ;
    LAYER M4 ;
    RECT 221.785 13.2 223.085 0 ;
    LAYER M4 ;
    RECT 226.425 13.2 227.425 0 ;
    LAYER M4 ;
    RECT 231.885 13.2 232.885 0 ;
    LAYER M4 ;
    RECT 236.225 13.2 237.525 0 ;
    LAYER M3 ;
    RECT 243.285 16.625 256.485 17.325 ;
    LAYER M3 ;
    RECT 243.285 24.875 256.485 25.575 ;
    LAYER M3 ;
    RECT 243.285 32.15 256.485 34.15 ;
    LAYER M3 ;
    RECT 243.285 37.82 256.485 38.36 ;
    LAYER M3 ;
    RECT 243.285 45.315 256.485 45.855 ;
    LAYER M3 ;
    RECT 243.285 55.92 256.485 56.72 ;
    LAYER M3 ;
    RECT 243.285 61.175 256.485 63.175 ;
    LAYER M3 ;
    RECT 243.285 65.705 256.485 68.705 ;
    LAYER M3 ;
    RECT 243.285 73.055 256.485 73.755 ;
    LAYER M3 ;
    RECT 243.285 76.705 256.485 77.405 ;
    LAYER M3 ;
    RECT 243.285 80.355 256.485 81.055 ;
    LAYER M3 ;
    RECT 243.285 84.005 256.485 84.705 ;
    LAYER M3 ;
    RECT 243.285 87.655 256.485 88.355 ;
    LAYER M3 ;
    RECT 243.285 91.305 256.485 92.005 ;
    LAYER M3 ;
    RECT 243.285 94.955 256.485 95.655 ;
    LAYER M3 ;
    RECT 243.285 98.605 256.485 99.305 ;
    LAYER M3 ;
    RECT 243.285 102.255 256.485 102.955 ;
    LAYER M3 ;
    RECT 243.285 105.905 256.485 106.605 ;
    LAYER M3 ;
    RECT 243.285 109.555 256.485 110.255 ;
    LAYER M3 ;
    RECT 243.285 113.205 256.485 113.905 ;
    LAYER M3 ;
    RECT 243.285 116.855 256.485 117.555 ;
    LAYER M3 ;
    RECT 243.285 120.505 256.485 121.205 ;
    LAYER M3 ;
    RECT 243.285 124.155 256.485 124.855 ;
    LAYER M3 ;
    RECT 243.285 127.805 256.485 128.505 ;
    LAYER M3 ;
    RECT 243.285 131.455 256.485 132.155 ;
    LAYER M3 ;
    RECT 243.285 135.105 256.485 135.805 ;
    LAYER M3 ;
    RECT 13.2 16.625 0 17.325 ;
    LAYER M3 ;
    RECT 13.2 24.875 0 25.575 ;
    LAYER M3 ;
    RECT 13.2 32.15 0 34.15 ;
    LAYER M3 ;
    RECT 13.2 37.82 0 38.36 ;
    LAYER M3 ;
    RECT 13.2 45.315 0 45.855 ;
    LAYER M3 ;
    RECT 13.2 55.92 0 56.72 ;
    LAYER M3 ;
    RECT 13.2 61.175 0 63.175 ;
    LAYER M3 ;
    RECT 13.2 65.705 0 68.705 ;
    LAYER M3 ;
    RECT 13.2 73.055 0 73.755 ;
    LAYER M3 ;
    RECT 13.2 76.705 0 77.405 ;
    LAYER M3 ;
    RECT 13.2 80.355 0 81.055 ;
    LAYER M3 ;
    RECT 13.2 84.005 0 84.705 ;
    LAYER M3 ;
    RECT 13.2 87.655 0 88.355 ;
    LAYER M3 ;
    RECT 13.2 91.305 0 92.005 ;
    LAYER M3 ;
    RECT 13.2 94.955 0 95.655 ;
    LAYER M3 ;
    RECT 13.2 98.605 0 99.305 ;
    LAYER M3 ;
    RECT 13.2 102.255 0 102.955 ;
    LAYER M3 ;
    RECT 13.2 105.905 0 106.605 ;
    LAYER M3 ;
    RECT 13.2 109.555 0 110.255 ;
    LAYER M3 ;
    RECT 13.2 113.205 0 113.905 ;
    LAYER M3 ;
    RECT 13.2 116.855 0 117.555 ;
    LAYER M3 ;
    RECT 13.2 120.505 0 121.205 ;
    LAYER M3 ;
    RECT 13.2 124.155 0 124.855 ;
    LAYER M3 ;
    RECT 13.2 127.805 0 128.505 ;
    LAYER M3 ;
    RECT 13.2 131.455 0 132.155 ;
    LAYER M3 ;
    RECT 13.2 135.105 0 135.805 ;
    LAYER M4 ;
    RECT 15.36 138.595 15.96 145.195 ;
    LAYER M4 ;
    RECT 16.445 138.595 17.265 145.195 ;
    LAYER M4 ;
    RECT 20.435 138.595 21.255 145.195 ;
    LAYER M4 ;
    RECT 21.765 138.595 22.585 145.195 ;
    LAYER M4 ;
    RECT 25.755 138.595 26.575 145.195 ;
    LAYER M4 ;
    RECT 27.085 138.595 27.905 145.195 ;
    LAYER M4 ;
    RECT 31.075 138.595 31.895 145.195 ;
    LAYER M4 ;
    RECT 32.405 138.595 33.225 145.195 ;
    LAYER M4 ;
    RECT 36.395 138.595 37.215 145.195 ;
    LAYER M4 ;
    RECT 37.725 138.595 38.545 145.195 ;
    LAYER M4 ;
    RECT 41.715 138.595 42.535 145.195 ;
    LAYER M4 ;
    RECT 43.045 138.595 43.865 145.195 ;
    LAYER M4 ;
    RECT 47.035 138.595 47.855 145.195 ;
    LAYER M4 ;
    RECT 48.365 138.595 49.185 145.195 ;
    LAYER M4 ;
    RECT 52.355 138.595 53.175 145.195 ;
    LAYER M4 ;
    RECT 53.685 138.595 54.505 145.195 ;
    LAYER M4 ;
    RECT 57.675 138.595 58.495 145.195 ;
    LAYER M4 ;
    RECT 58.98 138.595 59.58 145.195 ;
    LAYER M4 ;
    RECT 60.065 138.595 60.885 145.195 ;
    LAYER M4 ;
    RECT 64.055 138.595 64.875 145.195 ;
    LAYER M4 ;
    RECT 65.385 138.595 66.205 145.195 ;
    LAYER M4 ;
    RECT 69.375 138.595 70.195 145.195 ;
    LAYER M4 ;
    RECT 70.705 138.595 71.525 145.195 ;
    LAYER M4 ;
    RECT 74.695 138.595 75.515 145.195 ;
    LAYER M4 ;
    RECT 76.025 138.595 76.845 145.195 ;
    LAYER M4 ;
    RECT 80.015 138.595 80.835 145.195 ;
    LAYER M4 ;
    RECT 81.345 138.595 82.165 145.195 ;
    LAYER M4 ;
    RECT 85.335 138.595 86.155 145.195 ;
    LAYER M4 ;
    RECT 86.665 138.595 87.485 145.195 ;
    LAYER M4 ;
    RECT 90.655 138.595 91.475 145.195 ;
    LAYER M4 ;
    RECT 91.985 138.595 92.805 145.195 ;
    LAYER M4 ;
    RECT 95.975 138.595 96.795 145.195 ;
    LAYER M4 ;
    RECT 97.305 138.595 98.125 145.195 ;
    LAYER M4 ;
    RECT 101.295 138.595 102.115 145.195 ;
    LAYER M4 ;
    RECT 102.6 138.595 103.2 145.195 ;
    LAYER M4 ;
    RECT 107.33 138.595 108.39 145.195 ;
    LAYER M4 ;
    RECT 110.39 138.595 111.45 145.195 ;
    LAYER M4 ;
    RECT 113.45 138.595 114.51 145.195 ;
    LAYER M4 ;
    RECT 116.51 138.595 117.57 145.195 ;
    LAYER M4 ;
    RECT 119.57 138.595 120.63 145.195 ;
    LAYER M4 ;
    RECT 122.63 138.595 123.69 145.195 ;
    LAYER M4 ;
    RECT 125.69 138.595 126.75 145.195 ;
    LAYER M4 ;
    RECT 128.75 138.595 129.81 145.195 ;
    LAYER M4 ;
    RECT 131.81 138.595 132.87 145.195 ;
    LAYER M4 ;
    RECT 134.87 138.595 135.93 145.195 ;
    LAYER M4 ;
    RECT 137.93 138.595 138.99 145.195 ;
    LAYER M4 ;
    RECT 141.875 138.595 143.135 145.195 ;
    LAYER M4 ;
    RECT 145.955 138.595 147.215 145.195 ;
    LAYER M4 ;
    RECT 149.725 138.595 150.355 145.195 ;
    LAYER M4 ;
    RECT 150.895 138.595 151.495 145.195 ;
    LAYER M4 ;
    RECT 153.285 138.595 153.885 145.195 ;
    LAYER M4 ;
    RECT 154.37 138.595 155.19 145.195 ;
    LAYER M4 ;
    RECT 158.36 138.595 159.18 145.195 ;
    LAYER M4 ;
    RECT 159.69 138.595 160.51 145.195 ;
    LAYER M4 ;
    RECT 163.68 138.595 164.5 145.195 ;
    LAYER M4 ;
    RECT 165.01 138.595 165.83 145.195 ;
    LAYER M4 ;
    RECT 169 138.595 169.82 145.195 ;
    LAYER M4 ;
    RECT 170.33 138.595 171.15 145.195 ;
    LAYER M4 ;
    RECT 174.32 138.595 175.14 145.195 ;
    LAYER M4 ;
    RECT 175.65 138.595 176.47 145.195 ;
    LAYER M4 ;
    RECT 179.64 138.595 180.46 145.195 ;
    LAYER M4 ;
    RECT 180.97 138.595 181.79 145.195 ;
    LAYER M4 ;
    RECT 184.96 138.595 185.78 145.195 ;
    LAYER M4 ;
    RECT 186.29 138.595 187.11 145.195 ;
    LAYER M4 ;
    RECT 190.28 138.595 191.1 145.195 ;
    LAYER M4 ;
    RECT 191.61 138.595 192.43 145.195 ;
    LAYER M4 ;
    RECT 195.6 138.595 196.42 145.195 ;
    LAYER M4 ;
    RECT 196.905 138.595 197.505 145.195 ;
    LAYER M4 ;
    RECT 197.99 138.595 198.81 145.195 ;
    LAYER M4 ;
    RECT 201.98 138.595 202.8 145.195 ;
    LAYER M4 ;
    RECT 203.31 138.595 204.13 145.195 ;
    LAYER M4 ;
    RECT 207.3 138.595 208.12 145.195 ;
    LAYER M4 ;
    RECT 208.63 138.595 209.45 145.195 ;
    LAYER M4 ;
    RECT 212.62 138.595 213.44 145.195 ;
    LAYER M4 ;
    RECT 213.95 138.595 214.77 145.195 ;
    LAYER M4 ;
    RECT 217.94 138.595 218.76 145.195 ;
    LAYER M4 ;
    RECT 219.27 138.595 220.09 145.195 ;
    LAYER M4 ;
    RECT 223.26 138.595 224.08 145.195 ;
    LAYER M4 ;
    RECT 224.59 138.595 225.41 145.195 ;
    LAYER M4 ;
    RECT 228.58 138.595 229.4 145.195 ;
    LAYER M4 ;
    RECT 229.91 138.595 230.73 145.195 ;
    LAYER M4 ;
    RECT 233.9 138.595 234.72 145.195 ;
    LAYER M4 ;
    RECT 235.23 138.595 236.05 145.195 ;
    LAYER M4 ;
    RECT 239.22 138.595 240.04 145.195 ;
    LAYER M4 ;
    RECT 240.525 138.595 241.125 145.195 ;
    LAYER M4 ;
    RECT 14.19 13.2 14.79 6.6 ;
    LAYER M4 ;
    RECT 16.56 13.2 17.38 6.6 ;
    LAYER M4 ;
    RECT 20.72 13.2 22.02 6.6 ;
    LAYER M4 ;
    RECT 26.18 13.2 27.48 6.6 ;
    LAYER M4 ;
    RECT 31.64 13.2 32.94 6.6 ;
    LAYER M4 ;
    RECT 36.28 13.2 37.1 6.6 ;
    LAYER M4 ;
    RECT 37.84 13.2 38.66 6.6 ;
    LAYER M4 ;
    RECT 42 13.2 43.3 6.6 ;
    LAYER M4 ;
    RECT 47.46 13.2 48.76 6.6 ;
    LAYER M4 ;
    RECT 52.92 13.2 54.22 6.6 ;
    LAYER M4 ;
    RECT 57.56 13.2 58.38 6.6 ;
    LAYER M4 ;
    RECT 58.98 13.2 59.58 6.6 ;
    LAYER M4 ;
    RECT 60.18 13.2 61 6.6 ;
    LAYER M4 ;
    RECT 64.34 13.2 65.64 6.6 ;
    LAYER M4 ;
    RECT 69.8 13.2 71.1 6.6 ;
    LAYER M4 ;
    RECT 75.26 13.2 76.56 6.6 ;
    LAYER M4 ;
    RECT 79.9 13.2 80.72 6.6 ;
    LAYER M4 ;
    RECT 81.46 13.2 82.28 6.6 ;
    LAYER M4 ;
    RECT 85.62 13.2 86.92 6.6 ;
    LAYER M4 ;
    RECT 91.08 13.2 92.38 6.6 ;
    LAYER M4 ;
    RECT 96.54 13.2 97.84 6.6 ;
    LAYER M4 ;
    RECT 101.18 13.2 102 6.6 ;
    LAYER M4 ;
    RECT 104.93 13.2 106.19 6.6 ;
    LAYER M4 ;
    RECT 111.05 13.2 112.31 6.6 ;
    LAYER M4 ;
    RECT 117.17 13.2 118.43 6.6 ;
    LAYER M4 ;
    RECT 123.29 13.2 124.55 6.6 ;
    LAYER M4 ;
    RECT 129.41 13.2 130.67 6.6 ;
    LAYER M4 ;
    RECT 135.53 13.2 136.79 6.6 ;
    LAYER M4 ;
    RECT 141.915 13.2 142.735 6.6 ;
    LAYER M4 ;
    RECT 145.85 13.2 147.32 6.6 ;
    LAYER M4 ;
    RECT 150.36 13.2 151.36 6.6 ;
    LAYER M4 ;
    RECT 154.485 13.2 155.305 6.6 ;
    LAYER M4 ;
    RECT 158.645 13.2 159.945 6.6 ;
    LAYER M4 ;
    RECT 164.105 13.2 165.405 6.6 ;
    LAYER M4 ;
    RECT 169.565 13.2 170.865 6.6 ;
    LAYER M4 ;
    RECT 174.205 13.2 175.025 6.6 ;
    LAYER M4 ;
    RECT 175.765 13.2 176.585 6.6 ;
    LAYER M4 ;
    RECT 179.925 13.2 181.225 6.6 ;
    LAYER M4 ;
    RECT 185.385 13.2 186.685 6.6 ;
    LAYER M4 ;
    RECT 190.845 13.2 192.145 6.6 ;
    LAYER M4 ;
    RECT 195.485 13.2 196.305 6.6 ;
    LAYER M4 ;
    RECT 196.905 13.2 197.505 6.6 ;
    LAYER M4 ;
    RECT 198.105 13.2 198.925 6.6 ;
    LAYER M4 ;
    RECT 202.265 13.2 203.565 6.6 ;
    LAYER M4 ;
    RECT 207.725 13.2 209.025 6.6 ;
    LAYER M4 ;
    RECT 213.185 13.2 214.485 6.6 ;
    LAYER M4 ;
    RECT 217.825 13.2 218.645 6.6 ;
    LAYER M4 ;
    RECT 219.385 13.2 220.205 6.6 ;
    LAYER M4 ;
    RECT 223.545 13.2 224.845 6.6 ;
    LAYER M4 ;
    RECT 229.005 13.2 230.305 6.6 ;
    LAYER M4 ;
    RECT 234.465 13.2 235.765 6.6 ;
    LAYER M4 ;
    RECT 239.105 13.2 239.925 6.6 ;
    LAYER M4 ;
    RECT 241.695 13.2 242.295 6.6 ;
    LAYER M3 ;
    RECT 243.285 20.5 249.885 21.9 ;
    LAYER M3 ;
    RECT 243.285 27.605 249.885 29.605 ;
    LAYER M3 ;
    RECT 243.285 40.8 249.885 41.6 ;
    LAYER M3 ;
    RECT 243.285 47.94 249.885 48.74 ;
    LAYER M3 ;
    RECT 243.285 58.855 249.885 59.855 ;
    LAYER M3 ;
    RECT 243.285 74.88 249.885 75.58 ;
    LAYER M3 ;
    RECT 243.285 78.53 249.885 79.23 ;
    LAYER M3 ;
    RECT 243.285 82.18 249.885 82.88 ;
    LAYER M3 ;
    RECT 243.285 85.83 249.885 86.53 ;
    LAYER M3 ;
    RECT 243.285 89.48 249.885 90.18 ;
    LAYER M3 ;
    RECT 243.285 93.13 249.885 93.83 ;
    LAYER M3 ;
    RECT 243.285 96.78 249.885 97.48 ;
    LAYER M3 ;
    RECT 243.285 100.43 249.885 101.13 ;
    LAYER M3 ;
    RECT 243.285 104.08 249.885 104.78 ;
    LAYER M3 ;
    RECT 243.285 107.73 249.885 108.43 ;
    LAYER M3 ;
    RECT 243.285 111.38 249.885 112.08 ;
    LAYER M3 ;
    RECT 243.285 115.03 249.885 115.73 ;
    LAYER M3 ;
    RECT 243.285 118.68 249.885 119.38 ;
    LAYER M3 ;
    RECT 243.285 122.33 249.885 123.03 ;
    LAYER M3 ;
    RECT 243.285 125.98 249.885 126.68 ;
    LAYER M3 ;
    RECT 243.285 129.63 249.885 130.33 ;
    LAYER M3 ;
    RECT 243.285 133.28 249.885 133.98 ;
    LAYER M3 ;
    RECT 13.2 20.5 6.6 21.9 ;
    LAYER M3 ;
    RECT 13.2 27.605 6.6 29.605 ;
    LAYER M3 ;
    RECT 13.2 40.8 6.6 41.6 ;
    LAYER M3 ;
    RECT 13.2 47.94 6.6 48.74 ;
    LAYER M3 ;
    RECT 13.2 58.855 6.6 59.855 ;
    LAYER M3 ;
    RECT 13.2 74.88 6.6 75.58 ;
    LAYER M3 ;
    RECT 13.2 78.53 6.6 79.23 ;
    LAYER M3 ;
    RECT 13.2 82.18 6.6 82.88 ;
    LAYER M3 ;
    RECT 13.2 85.83 6.6 86.53 ;
    LAYER M3 ;
    RECT 13.2 89.48 6.6 90.18 ;
    LAYER M3 ;
    RECT 13.2 93.13 6.6 93.83 ;
    LAYER M3 ;
    RECT 13.2 96.78 6.6 97.48 ;
    LAYER M3 ;
    RECT 13.2 100.43 6.6 101.13 ;
    LAYER M3 ;
    RECT 13.2 104.08 6.6 104.78 ;
    LAYER M3 ;
    RECT 13.2 107.73 6.6 108.43 ;
    LAYER M3 ;
    RECT 13.2 111.38 6.6 112.08 ;
    LAYER M3 ;
    RECT 13.2 115.03 6.6 115.73 ;
    LAYER M3 ;
    RECT 13.2 118.68 6.6 119.38 ;
    LAYER M3 ;
    RECT 13.2 122.33 6.6 123.03 ;
    LAYER M3 ;
    RECT 13.2 125.98 6.6 126.68 ;
    LAYER M3 ;
    RECT 13.2 129.63 6.6 130.33 ;
    LAYER M3 ;
    RECT 13.2 133.28 6.6 133.98 ;
    END
  END ram_256x16A
END LIBRARY

